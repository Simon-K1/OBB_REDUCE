// Generator : SpinalHDL v1.7.3    git head : ed8004c489ee8a38c2cab309d0447b543fe9d5b8
// Component : Conv

`timescale 1ns/1ps

module Conv (
  input               sData_valid,
  output reg          sData_ready,
  input      [127:0]  sData_payload,
  input               sFeatureFirstLayerData_valid,
  output              sFeatureFirstLayerData_ready,
  input      [7:0]    sFeatureFirstLayerData_payload,
  output              mData_valid,
  input               mData_ready,
  output     [127:0]  mData_payload,
  input      [31:0]   instruction_0,
  input      [31:0]   instruction_1,
  input      [31:0]   instruction_2,
  input      [31:0]   instruction_3,
  input      [31:0]   instruction_4,
  input      [3:0]    control,
  output     [3:0]    state,
  output              dmaReadValid,
  output              dmaFirstLayerReadValid,
  output              dmaWriteValid,
  input               introut,
  output              last,
  input               reset,
  input               clk
);

  reg        [3:0]    convState_1_complete;
  reg                 convCompute_1_sParaData_valid;
  reg        [127:0]  convCompute_1_sParaData_payload;
  reg                 convCompute_1_sFeatureData_valid;
  reg        [127:0]  convCompute_1_sFeatureData_payload;
  wire       [9:0]    convCompute_1_rowNumIn;
  wire       [9:0]    convCompute_1_colNumIn;
  wire       [11:0]   convCompute_1_channelIn;
  wire       [11:0]   convCompute_1_channelOut;
  wire                convCompute_1_enPadding;
  wire                convCompute_1_enActivation;
  wire       [7:0]    convCompute_1_zeroDara;
  wire       [0:0]    convCompute_1_zeroNum;
  wire       [12:0]   convCompute_1_weightNum;
  wire       [7:0]    convCompute_1_quanNum;
  wire       [7:0]    convCompute_1_quanZeroData;
  wire                convCompute_1_enStride;
  wire                convCompute_1_firstLayer;
  wire       [1:0]    convCompute_1_convType;
  wire       [31:0]   convCompute_1_amendReg;
  wire       [3:0]    convState_1_state;
  wire       [3:0]    convState_1_sign;
  wire                convState_1_dmaReadValid;
  wire                convState_1_dmaWriteValid;
  wire                convState_1_softReset;
  wire                convCompute_1_sParaData_ready;
  wire                convCompute_1_sFeatureData_ready;
  wire                convCompute_1_sFeatureFirstLayerData_ready;
  wire                convCompute_1_mFeatureData_valid;
  wire       [127:0]  convCompute_1_mFeatureData_payload;
  wire                convCompute_1_copyWeightDone;
  wire                convCompute_1_computeComplete;
  wire                convCompute_1_last;
  wire       [10:0]   _zz_channelIn;
  wire       [9:0]    _zz_channelOut;
  wire       [10:0]   _zz_rowNumIn;
  wire       [2:0]    _zz_zeroNum;
  wire       [15:0]   _zz_weightNum;
  wire       [15:0]   _zz_quanNum;
  reg                 para;
  wire                when_Conv_l33;
  wire                when_Conv_l33_1;
  reg                 compute;
  wire                when_Conv_l34;
  wire                when_Conv_l34_1;
  wire       [159:0]  computeInstruction;
  reg        [159:0]  computeInstructionReg;
  reg                 convState_1_softReset_delay_1;
  reg                 convState_1_softReset_delay_2;
  reg                 para_delay_1;
  reg                 para_delay_2;
  reg                 para_delay_3;
  reg                 compute_delay_1;
  reg                 compute_delay_2;
  reg                 compute_delay_3;
  reg                 writeComplete;
  wire                when_Conv_l89;
  reg                 computeComplete;
  wire                when_Conv_l93;
  wire                when_Conv_l97;
  (* max_fanout = "10" *) reg        [1:0]    dest;
  wire                when_Conv_l104;
  wire                when_Conv_l106;
  wire                when_Conv_l112;
  wire                when_Conv_l117;

  assign _zz_channelIn = computeInstructionReg[31 : 21];
  assign _zz_channelOut = computeInstructionReg[41 : 32];
  assign _zz_rowNumIn = computeInstructionReg[10 : 0];
  assign _zz_zeroNum = computeInstructionReg[54 : 52];
  assign _zz_weightNum = computeInstructionReg[111 : 96];
  assign _zz_quanNum = computeInstructionReg[127 : 112];
  ConvState convState_1 (
    .control       (control[3:0]             ), //i
    .complete      (convState_1_complete[3:0]), //i
    .state         (convState_1_state[3:0]   ), //o
    .sign          (convState_1_sign[3:0]    ), //o
    .dmaReadValid  (convState_1_dmaReadValid ), //o
    .dmaWriteValid (convState_1_dmaWriteValid), //o
    .softReset     (convState_1_softReset    ), //o
    .clk           (clk                      ), //i
    .reset         (reset                    )  //i
  );
  ConvCompute convCompute_1 (
    .startPa                        (para_delay_3                              ), //i
    .startCu                        (compute_delay_3                           ), //i
    .sParaData_valid                (convCompute_1_sParaData_valid             ), //i
    .sParaData_ready                (convCompute_1_sParaData_ready             ), //o
    .sParaData_payload              (convCompute_1_sParaData_payload[127:0]    ), //i
    .sFeatureData_valid             (convCompute_1_sFeatureData_valid          ), //i
    .sFeatureData_ready             (convCompute_1_sFeatureData_ready          ), //o
    .sFeatureData_payload           (convCompute_1_sFeatureData_payload[127:0] ), //i
    .sFeatureFirstLayerData_valid   (sFeatureFirstLayerData_valid              ), //i
    .sFeatureFirstLayerData_ready   (convCompute_1_sFeatureFirstLayerData_ready), //o
    .sFeatureFirstLayerData_payload (sFeatureFirstLayerData_payload[7:0]       ), //i
    .mFeatureData_valid             (convCompute_1_mFeatureData_valid          ), //o
    .mFeatureData_ready             (mData_ready                               ), //i
    .mFeatureData_payload           (convCompute_1_mFeatureData_payload[127:0] ), //o
    .copyWeightDone                 (convCompute_1_copyWeightDone              ), //o
    .computeComplete                (convCompute_1_computeComplete             ), //o
    .rowNumIn                       (convCompute_1_rowNumIn[9:0]               ), //i
    .colNumIn                       (convCompute_1_colNumIn[9:0]               ), //i
    .channelIn                      (convCompute_1_channelIn[11:0]             ), //i
    .channelOut                     (convCompute_1_channelOut[11:0]            ), //i
    .enPadding                      (convCompute_1_enPadding                   ), //i
    .enActivation                   (convCompute_1_enActivation                ), //i
    .zeroDara                       (convCompute_1_zeroDara[7:0]               ), //i
    .zeroNum                        (convCompute_1_zeroNum                     ), //i
    .weightNum                      (convCompute_1_weightNum[12:0]             ), //i
    .quanNum                        (convCompute_1_quanNum[7:0]                ), //i
    .quanZeroData                   (convCompute_1_quanZeroData[7:0]           ), //i
    .enStride                       (convCompute_1_enStride                    ), //i
    .firstLayer                     (convCompute_1_firstLayer                  ), //i
    .convType                       (convCompute_1_convType[1:0]               ), //i
    .last                           (convCompute_1_last                        ), //o
    .softReset                      (convState_1_softReset_delay_2             ), //i
    .amendReg                       (convCompute_1_amendReg[31:0]              ), //i
    .reset                          (reset                                     ), //i
    .clk                            (clk                                       )  //i
  );
  assign state = convState_1_state;
  assign when_Conv_l33 = (convState_1_sign == 4'b0001);
  assign when_Conv_l33_1 = (convState_1_sign != 4'b0001);
  assign when_Conv_l34 = (convState_1_sign == 4'b0010);
  assign when_Conv_l34_1 = (convState_1_sign != 4'b0010);
  assign computeInstruction = {instruction_4,{instruction_3,{instruction_2,{instruction_1,instruction_0}}}};
  assign last = convCompute_1_last;
  assign sFeatureFirstLayerData_ready = convCompute_1_sFeatureFirstLayerData_ready;
  assign convCompute_1_channelIn = {1'd0, _zz_channelIn};
  assign convCompute_1_channelOut = {2'd0, _zz_channelOut};
  assign convCompute_1_rowNumIn = _zz_rowNumIn[9:0];
  assign convCompute_1_colNumIn = computeInstructionReg[20 : 11];
  assign convCompute_1_enPadding = computeInstructionReg[42];
  assign convCompute_1_enActivation = computeInstructionReg[43];
  assign convCompute_1_zeroDara = computeInstructionReg[51 : 44];
  assign convCompute_1_zeroNum = _zz_zeroNum[0:0];
  assign convCompute_1_quanZeroData = computeInstructionReg[62 : 55];
  assign convCompute_1_convType = computeInstructionReg[65 : 64];
  assign convCompute_1_enStride = computeInstructionReg[63];
  assign convCompute_1_firstLayer = computeInstructionReg[66];
  assign convCompute_1_amendReg = computeInstructionReg[159 : 128];
  assign convCompute_1_weightNum = _zz_weightNum[12:0];
  assign convCompute_1_quanNum = _zz_quanNum[7:0];
  assign dmaReadValid = (convState_1_dmaReadValid && (! computeInstructionReg[66]));
  assign dmaFirstLayerReadValid = (convState_1_dmaReadValid && computeInstructionReg[66]);
  assign dmaWriteValid = convState_1_dmaWriteValid;
  assign when_Conv_l89 = (control == 4'b1111);
  assign when_Conv_l93 = (control == 4'b1111);
  always @(*) begin
    if(convCompute_1_copyWeightDone) begin
      convState_1_complete = 4'b0001;
    end else begin
      if(when_Conv_l97) begin
        convState_1_complete = 4'b0010;
      end else begin
        convState_1_complete = 4'b0000;
      end
    end
  end

  assign when_Conv_l97 = (computeComplete && writeComplete);
  assign when_Conv_l104 = (control == 4'b0001);
  assign when_Conv_l106 = (control == 4'b0010);
  assign when_Conv_l112 = (dest == 2'b00);
  always @(*) begin
    if(when_Conv_l112) begin
      convCompute_1_sParaData_valid = sData_valid;
    end else begin
      if(when_Conv_l117) begin
        convCompute_1_sParaData_valid = 1'b0;
      end else begin
        convCompute_1_sParaData_valid = 1'b0;
      end
    end
  end

  always @(*) begin
    if(when_Conv_l112) begin
      sData_ready = convCompute_1_sParaData_ready;
    end else begin
      if(when_Conv_l117) begin
        sData_ready = convCompute_1_sFeatureData_ready;
      end else begin
        sData_ready = 1'b0;
      end
    end
  end

  always @(*) begin
    if(when_Conv_l112) begin
      convCompute_1_sParaData_payload = sData_payload;
    end else begin
      if(when_Conv_l117) begin
        convCompute_1_sParaData_payload = 128'h0;
      end else begin
        convCompute_1_sParaData_payload = 128'h0;
      end
    end
  end

  always @(*) begin
    if(when_Conv_l112) begin
      convCompute_1_sFeatureData_valid = 1'b0;
    end else begin
      if(when_Conv_l117) begin
        convCompute_1_sFeatureData_valid = sData_valid;
      end else begin
        convCompute_1_sFeatureData_valid = 1'b0;
      end
    end
  end

  always @(*) begin
    if(when_Conv_l112) begin
      convCompute_1_sFeatureData_payload = 128'h0;
    end else begin
      if(when_Conv_l117) begin
        convCompute_1_sFeatureData_payload = sData_payload;
      end else begin
        convCompute_1_sFeatureData_payload = 128'h0;
      end
    end
  end

  assign when_Conv_l117 = (dest == 2'b01);
  assign mData_valid = convCompute_1_mFeatureData_valid;
  assign mData_payload = convCompute_1_mFeatureData_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      para <= 1'b0;
      compute <= 1'b0;
      computeInstructionReg <= 160'h0;
      writeComplete <= 1'b0;
      computeComplete <= 1'b0;
      dest <= 2'b11;
    end else begin
      if(when_Conv_l33) begin
        para <= 1'b1;
      end
      if(when_Conv_l33_1) begin
        para <= 1'b0;
      end
      if(when_Conv_l34) begin
        compute <= 1'b1;
      end
      if(when_Conv_l34_1) begin
        compute <= 1'b0;
      end
      computeInstructionReg <= computeInstruction;
      if(introut) begin
        writeComplete <= 1'b1;
      end
      if(when_Conv_l89) begin
        writeComplete <= 1'b0;
      end
      if(convCompute_1_computeComplete) begin
        computeComplete <= 1'b1;
      end
      if(when_Conv_l93) begin
        computeComplete <= 1'b0;
      end
      if(when_Conv_l104) begin
        dest <= 2'b00;
      end else begin
        if(when_Conv_l106) begin
          dest <= 2'b01;
        end else begin
          dest <= dest;
        end
      end
    end
  end

  always @(posedge clk) begin
    convState_1_softReset_delay_1 <= convState_1_softReset;
    convState_1_softReset_delay_2 <= convState_1_softReset_delay_1;
    para_delay_1 <= para;
    para_delay_2 <= para_delay_1;
    para_delay_3 <= para_delay_2;
    compute_delay_1 <= compute;
    compute_delay_2 <= compute_delay_1;
    compute_delay_3 <= compute_delay_2;
  end


endmodule

module ConvCompute (
  input               startPa,
  input               startCu,
  input               sParaData_valid,
  output              sParaData_ready,
  input      [127:0]  sParaData_payload,
  input               sFeatureData_valid,
  output reg          sFeatureData_ready,
  input      [127:0]  sFeatureData_payload,
  input               sFeatureFirstLayerData_valid,
  output              sFeatureFirstLayerData_ready,
  input      [7:0]    sFeatureFirstLayerData_payload,
  output              mFeatureData_valid,
  input               mFeatureData_ready,
  output     [127:0]  mFeatureData_payload,
  output              copyWeightDone,
  output              computeComplete,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input      [11:0]   channelIn,
  input      [11:0]   channelOut,
  input               enPadding,
  input               enActivation,
  input      [7:0]    zeroDara,
  input      [0:0]    zeroNum,
  input      [12:0]   weightNum,
  input      [7:0]    quanNum,
  input      [7:0]    quanZeroData,
  input               enStride,
  input               firstLayer,
  input      [1:0]    convType,
  output              last,
  input               softReset,
  input      [31:0]   amendReg,
  input               reset,
  input               clk
);

  reg                 channelIncr_1_mData_ready;
  reg                 dataGenerate_1_sData_valid;
  reg        [127:0]  dataGenerate_1_sData_payload;
  wire       [13:0]   waXpmSyncFifo_9_sCount;
  wire       [13:0]   waXpmSyncFifo_9_mCount;
  wire       [7:0]    dSP_1_a;
  wire       [7:0]    dSP_1_d;
  wire       [7:0]    dSP_1_b;
  wire       [7:0]    dSP_2_a;
  wire       [7:0]    dSP_2_d;
  wire       [7:0]    dSP_2_b;
  wire       [7:0]    dSP_3_a;
  wire       [7:0]    dSP_3_d;
  wire       [7:0]    dSP_3_b;
  wire       [7:0]    dSP_4_a;
  wire       [7:0]    dSP_4_d;
  wire       [7:0]    dSP_4_b;
  wire       [7:0]    dSP_5_a;
  wire       [7:0]    dSP_5_d;
  wire       [7:0]    dSP_5_b;
  wire       [7:0]    dSP_6_a;
  wire       [7:0]    dSP_6_d;
  wire       [7:0]    dSP_6_b;
  wire       [7:0]    dSP_7_a;
  wire       [7:0]    dSP_7_d;
  wire       [7:0]    dSP_7_b;
  wire       [7:0]    dSP_8_a;
  wire       [7:0]    dSP_8_d;
  wire       [7:0]    dSP_8_b;
  wire       [7:0]    dSP_9_a;
  wire       [7:0]    dSP_9_d;
  wire       [7:0]    dSP_9_b;
  wire       [7:0]    dSP_10_a;
  wire       [7:0]    dSP_10_d;
  wire       [7:0]    dSP_10_b;
  wire       [7:0]    dSP_11_a;
  wire       [7:0]    dSP_11_d;
  wire       [7:0]    dSP_11_b;
  wire       [7:0]    dSP_12_a;
  wire       [7:0]    dSP_12_d;
  wire       [7:0]    dSP_12_b;
  wire       [7:0]    dSP_13_a;
  wire       [7:0]    dSP_13_d;
  wire       [7:0]    dSP_13_b;
  wire       [7:0]    dSP_14_a;
  wire       [7:0]    dSP_14_d;
  wire       [7:0]    dSP_14_b;
  wire       [7:0]    dSP_15_a;
  wire       [7:0]    dSP_15_d;
  wire       [7:0]    dSP_15_b;
  wire       [7:0]    dSP_16_a;
  wire       [7:0]    dSP_16_d;
  wire       [7:0]    dSP_16_b;
  wire       [7:0]    dSP_17_a;
  wire       [7:0]    dSP_17_d;
  wire       [7:0]    dSP_17_b;
  wire       [7:0]    dSP_18_a;
  wire       [7:0]    dSP_18_d;
  wire       [7:0]    dSP_18_b;
  wire       [7:0]    dSP_19_a;
  wire       [7:0]    dSP_19_d;
  wire       [7:0]    dSP_19_b;
  wire       [7:0]    dSP_20_a;
  wire       [7:0]    dSP_20_d;
  wire       [7:0]    dSP_20_b;
  wire       [7:0]    dSP_21_a;
  wire       [7:0]    dSP_21_d;
  wire       [7:0]    dSP_21_b;
  wire       [7:0]    dSP_22_a;
  wire       [7:0]    dSP_22_d;
  wire       [7:0]    dSP_22_b;
  wire       [7:0]    dSP_23_a;
  wire       [7:0]    dSP_23_d;
  wire       [7:0]    dSP_23_b;
  wire       [7:0]    dSP_24_a;
  wire       [7:0]    dSP_24_d;
  wire       [7:0]    dSP_24_b;
  wire       [7:0]    dSP_25_a;
  wire       [7:0]    dSP_25_d;
  wire       [7:0]    dSP_25_b;
  wire       [7:0]    dSP_26_a;
  wire       [7:0]    dSP_26_d;
  wire       [7:0]    dSP_26_b;
  wire       [7:0]    dSP_27_a;
  wire       [7:0]    dSP_27_d;
  wire       [7:0]    dSP_27_b;
  wire       [7:0]    dSP_28_a;
  wire       [7:0]    dSP_28_d;
  wire       [7:0]    dSP_28_b;
  wire       [7:0]    dSP_29_a;
  wire       [7:0]    dSP_29_d;
  wire       [7:0]    dSP_29_b;
  wire       [7:0]    dSP_30_a;
  wire       [7:0]    dSP_30_d;
  wire       [7:0]    dSP_30_b;
  wire       [7:0]    dSP_31_a;
  wire       [7:0]    dSP_31_d;
  wire       [7:0]    dSP_31_b;
  wire       [7:0]    dSP_32_a;
  wire       [7:0]    dSP_32_d;
  wire       [7:0]    dSP_32_b;
  wire       [7:0]    dSP_33_a;
  wire       [7:0]    dSP_33_d;
  wire       [7:0]    dSP_33_b;
  wire       [7:0]    dSP_34_a;
  wire       [7:0]    dSP_34_d;
  wire       [7:0]    dSP_34_b;
  wire       [7:0]    dSP_35_a;
  wire       [7:0]    dSP_35_d;
  wire       [7:0]    dSP_35_b;
  wire       [7:0]    dSP_36_a;
  wire       [7:0]    dSP_36_d;
  wire       [7:0]    dSP_36_b;
  wire       [7:0]    dSP_37_a;
  wire       [7:0]    dSP_37_d;
  wire       [7:0]    dSP_37_b;
  wire       [7:0]    dSP_38_a;
  wire       [7:0]    dSP_38_d;
  wire       [7:0]    dSP_38_b;
  wire       [7:0]    dSP_39_a;
  wire       [7:0]    dSP_39_d;
  wire       [7:0]    dSP_39_b;
  wire       [7:0]    dSP_40_a;
  wire       [7:0]    dSP_40_d;
  wire       [7:0]    dSP_40_b;
  wire       [7:0]    dSP_41_a;
  wire       [7:0]    dSP_41_d;
  wire       [7:0]    dSP_41_b;
  wire       [7:0]    dSP_42_a;
  wire       [7:0]    dSP_42_d;
  wire       [7:0]    dSP_42_b;
  wire       [7:0]    dSP_43_a;
  wire       [7:0]    dSP_43_d;
  wire       [7:0]    dSP_43_b;
  wire       [7:0]    dSP_44_a;
  wire       [7:0]    dSP_44_d;
  wire       [7:0]    dSP_44_b;
  wire       [7:0]    dSP_45_a;
  wire       [7:0]    dSP_45_d;
  wire       [7:0]    dSP_45_b;
  wire       [7:0]    dSP_46_a;
  wire       [7:0]    dSP_46_d;
  wire       [7:0]    dSP_46_b;
  wire       [7:0]    dSP_47_a;
  wire       [7:0]    dSP_47_d;
  wire       [7:0]    dSP_47_b;
  wire       [7:0]    dSP_48_a;
  wire       [7:0]    dSP_48_d;
  wire       [7:0]    dSP_48_b;
  wire       [7:0]    dSP_49_a;
  wire       [7:0]    dSP_49_d;
  wire       [7:0]    dSP_49_b;
  wire       [7:0]    dSP_50_a;
  wire       [7:0]    dSP_50_d;
  wire       [7:0]    dSP_50_b;
  wire       [7:0]    dSP_51_a;
  wire       [7:0]    dSP_51_d;
  wire       [7:0]    dSP_51_b;
  wire       [7:0]    dSP_52_a;
  wire       [7:0]    dSP_52_d;
  wire       [7:0]    dSP_52_b;
  wire       [7:0]    dSP_53_a;
  wire       [7:0]    dSP_53_d;
  wire       [7:0]    dSP_53_b;
  wire       [7:0]    dSP_54_a;
  wire       [7:0]    dSP_54_d;
  wire       [7:0]    dSP_54_b;
  wire       [7:0]    dSP_55_a;
  wire       [7:0]    dSP_55_d;
  wire       [7:0]    dSP_55_b;
  wire       [7:0]    dSP_56_a;
  wire       [7:0]    dSP_56_d;
  wire       [7:0]    dSP_56_b;
  wire       [7:0]    dSP_57_a;
  wire       [7:0]    dSP_57_d;
  wire       [7:0]    dSP_57_b;
  wire       [7:0]    dSP_58_a;
  wire       [7:0]    dSP_58_d;
  wire       [7:0]    dSP_58_b;
  wire       [7:0]    dSP_59_a;
  wire       [7:0]    dSP_59_d;
  wire       [7:0]    dSP_59_b;
  wire       [7:0]    dSP_60_a;
  wire       [7:0]    dSP_60_d;
  wire       [7:0]    dSP_60_b;
  wire       [7:0]    dSP_61_a;
  wire       [7:0]    dSP_61_d;
  wire       [7:0]    dSP_61_b;
  wire       [7:0]    dSP_62_a;
  wire       [7:0]    dSP_62_d;
  wire       [7:0]    dSP_62_b;
  wire       [7:0]    dSP_63_a;
  wire       [7:0]    dSP_63_d;
  wire       [7:0]    dSP_63_b;
  wire       [7:0]    dSP_64_a;
  wire       [7:0]    dSP_64_d;
  wire       [7:0]    dSP_64_b;
  wire       [7:0]    dSP_65_a;
  wire       [7:0]    dSP_65_d;
  wire       [7:0]    dSP_65_b;
  wire       [7:0]    dSP_66_a;
  wire       [7:0]    dSP_66_d;
  wire       [7:0]    dSP_66_b;
  wire       [7:0]    dSP_67_a;
  wire       [7:0]    dSP_67_d;
  wire       [7:0]    dSP_67_b;
  wire       [7:0]    dSP_68_a;
  wire       [7:0]    dSP_68_d;
  wire       [7:0]    dSP_68_b;
  wire       [7:0]    dSP_69_a;
  wire       [7:0]    dSP_69_d;
  wire       [7:0]    dSP_69_b;
  wire       [7:0]    dSP_70_a;
  wire       [7:0]    dSP_70_d;
  wire       [7:0]    dSP_70_b;
  wire       [7:0]    dSP_71_a;
  wire       [7:0]    dSP_71_d;
  wire       [7:0]    dSP_71_b;
  wire       [7:0]    dSP_72_a;
  wire       [7:0]    dSP_72_d;
  wire       [7:0]    dSP_72_b;
  wire       [7:0]    dSP_73_a;
  wire       [7:0]    dSP_73_d;
  wire       [7:0]    dSP_73_b;
  wire       [7:0]    dSP_74_a;
  wire       [7:0]    dSP_74_d;
  wire       [7:0]    dSP_74_b;
  wire       [7:0]    dSP_75_a;
  wire       [7:0]    dSP_75_d;
  wire       [7:0]    dSP_75_b;
  wire       [7:0]    dSP_76_a;
  wire       [7:0]    dSP_76_d;
  wire       [7:0]    dSP_76_b;
  wire       [7:0]    dSP_77_a;
  wire       [7:0]    dSP_77_d;
  wire       [7:0]    dSP_77_b;
  wire       [7:0]    dSP_78_a;
  wire       [7:0]    dSP_78_d;
  wire       [7:0]    dSP_78_b;
  wire       [7:0]    dSP_79_a;
  wire       [7:0]    dSP_79_d;
  wire       [7:0]    dSP_79_b;
  wire       [7:0]    dSP_80_a;
  wire       [7:0]    dSP_80_d;
  wire       [7:0]    dSP_80_b;
  wire       [7:0]    dSP_81_a;
  wire       [7:0]    dSP_81_d;
  wire       [7:0]    dSP_81_b;
  wire       [7:0]    dSP_82_a;
  wire       [7:0]    dSP_82_d;
  wire       [7:0]    dSP_82_b;
  wire       [7:0]    dSP_83_a;
  wire       [7:0]    dSP_83_d;
  wire       [7:0]    dSP_83_b;
  wire       [7:0]    dSP_84_a;
  wire       [7:0]    dSP_84_d;
  wire       [7:0]    dSP_84_b;
  wire       [7:0]    dSP_85_a;
  wire       [7:0]    dSP_85_d;
  wire       [7:0]    dSP_85_b;
  wire       [7:0]    dSP_86_a;
  wire       [7:0]    dSP_86_d;
  wire       [7:0]    dSP_86_b;
  wire       [7:0]    dSP_87_a;
  wire       [7:0]    dSP_87_d;
  wire       [7:0]    dSP_87_b;
  wire       [7:0]    dSP_88_a;
  wire       [7:0]    dSP_88_d;
  wire       [7:0]    dSP_88_b;
  wire       [7:0]    dSP_89_a;
  wire       [7:0]    dSP_89_d;
  wire       [7:0]    dSP_89_b;
  wire       [7:0]    dSP_90_a;
  wire       [7:0]    dSP_90_d;
  wire       [7:0]    dSP_90_b;
  wire       [7:0]    dSP_91_a;
  wire       [7:0]    dSP_91_d;
  wire       [7:0]    dSP_91_b;
  wire       [7:0]    dSP_92_a;
  wire       [7:0]    dSP_92_d;
  wire       [7:0]    dSP_92_b;
  wire       [7:0]    dSP_93_a;
  wire       [7:0]    dSP_93_d;
  wire       [7:0]    dSP_93_b;
  wire       [7:0]    dSP_94_a;
  wire       [7:0]    dSP_94_d;
  wire       [7:0]    dSP_94_b;
  wire       [7:0]    dSP_95_a;
  wire       [7:0]    dSP_95_d;
  wire       [7:0]    dSP_95_b;
  wire       [7:0]    dSP_96_a;
  wire       [7:0]    dSP_96_d;
  wire       [7:0]    dSP_96_b;
  wire       [7:0]    dSP_97_a;
  wire       [7:0]    dSP_97_d;
  wire       [7:0]    dSP_97_b;
  wire       [7:0]    dSP_98_a;
  wire       [7:0]    dSP_98_d;
  wire       [7:0]    dSP_98_b;
  wire       [7:0]    dSP_99_a;
  wire       [7:0]    dSP_99_d;
  wire       [7:0]    dSP_99_b;
  wire       [7:0]    dSP_100_a;
  wire       [7:0]    dSP_100_d;
  wire       [7:0]    dSP_100_b;
  wire       [7:0]    dSP_101_a;
  wire       [7:0]    dSP_101_d;
  wire       [7:0]    dSP_101_b;
  wire       [7:0]    dSP_102_a;
  wire       [7:0]    dSP_102_d;
  wire       [7:0]    dSP_102_b;
  wire       [7:0]    dSP_103_a;
  wire       [7:0]    dSP_103_d;
  wire       [7:0]    dSP_103_b;
  wire       [7:0]    dSP_104_a;
  wire       [7:0]    dSP_104_d;
  wire       [7:0]    dSP_104_b;
  wire       [7:0]    dSP_105_a;
  wire       [7:0]    dSP_105_d;
  wire       [7:0]    dSP_105_b;
  wire       [7:0]    dSP_106_a;
  wire       [7:0]    dSP_106_d;
  wire       [7:0]    dSP_106_b;
  wire       [7:0]    dSP_107_a;
  wire       [7:0]    dSP_107_d;
  wire       [7:0]    dSP_107_b;
  wire       [7:0]    dSP_108_a;
  wire       [7:0]    dSP_108_d;
  wire       [7:0]    dSP_108_b;
  wire       [7:0]    dSP_109_a;
  wire       [7:0]    dSP_109_d;
  wire       [7:0]    dSP_109_b;
  wire       [7:0]    dSP_110_a;
  wire       [7:0]    dSP_110_d;
  wire       [7:0]    dSP_110_b;
  wire       [7:0]    dSP_111_a;
  wire       [7:0]    dSP_111_d;
  wire       [7:0]    dSP_111_b;
  wire       [7:0]    dSP_112_a;
  wire       [7:0]    dSP_112_d;
  wire       [7:0]    dSP_112_b;
  wire       [7:0]    dSP_113_a;
  wire       [7:0]    dSP_113_d;
  wire       [7:0]    dSP_113_b;
  wire       [7:0]    dSP_114_a;
  wire       [7:0]    dSP_114_d;
  wire       [7:0]    dSP_114_b;
  wire       [7:0]    dSP_115_a;
  wire       [7:0]    dSP_115_d;
  wire       [7:0]    dSP_115_b;
  wire       [7:0]    dSP_116_a;
  wire       [7:0]    dSP_116_d;
  wire       [7:0]    dSP_116_b;
  wire       [7:0]    dSP_117_a;
  wire       [7:0]    dSP_117_d;
  wire       [7:0]    dSP_117_b;
  wire       [7:0]    dSP_118_a;
  wire       [7:0]    dSP_118_d;
  wire       [7:0]    dSP_118_b;
  wire       [7:0]    dSP_119_a;
  wire       [7:0]    dSP_119_d;
  wire       [7:0]    dSP_119_b;
  wire       [7:0]    dSP_120_a;
  wire       [7:0]    dSP_120_d;
  wire       [7:0]    dSP_120_b;
  wire       [7:0]    dSP_121_a;
  wire       [7:0]    dSP_121_d;
  wire       [7:0]    dSP_121_b;
  wire       [7:0]    dSP_122_a;
  wire       [7:0]    dSP_122_d;
  wire       [7:0]    dSP_122_b;
  wire       [7:0]    dSP_123_a;
  wire       [7:0]    dSP_123_d;
  wire       [7:0]    dSP_123_b;
  wire       [7:0]    dSP_124_a;
  wire       [7:0]    dSP_124_d;
  wire       [7:0]    dSP_124_b;
  wire       [7:0]    dSP_125_a;
  wire       [7:0]    dSP_125_d;
  wire       [7:0]    dSP_125_b;
  wire       [7:0]    dSP_126_a;
  wire       [7:0]    dSP_126_d;
  wire       [7:0]    dSP_126_b;
  wire       [7:0]    dSP_127_a;
  wire       [7:0]    dSP_127_d;
  wire       [7:0]    dSP_127_b;
  wire       [7:0]    dSP_128_a;
  wire       [7:0]    dSP_128_d;
  wire       [7:0]    dSP_128_b;
  wire       [7:0]    dSP_129_a;
  wire       [7:0]    dSP_129_d;
  wire       [7:0]    dSP_129_b;
  wire       [7:0]    dSP_130_a;
  wire       [7:0]    dSP_130_d;
  wire       [7:0]    dSP_130_b;
  wire       [7:0]    dSP_131_a;
  wire       [7:0]    dSP_131_d;
  wire       [7:0]    dSP_131_b;
  wire       [7:0]    dSP_132_a;
  wire       [7:0]    dSP_132_d;
  wire       [7:0]    dSP_132_b;
  wire       [7:0]    dSP_133_a;
  wire       [7:0]    dSP_133_d;
  wire       [7:0]    dSP_133_b;
  wire       [7:0]    dSP_134_a;
  wire       [7:0]    dSP_134_d;
  wire       [7:0]    dSP_134_b;
  wire       [7:0]    dSP_135_a;
  wire       [7:0]    dSP_135_d;
  wire       [7:0]    dSP_135_b;
  wire       [7:0]    dSP_136_a;
  wire       [7:0]    dSP_136_d;
  wire       [7:0]    dSP_136_b;
  wire       [7:0]    dSP_137_a;
  wire       [7:0]    dSP_137_d;
  wire       [7:0]    dSP_137_b;
  wire       [7:0]    dSP_138_a;
  wire       [7:0]    dSP_138_d;
  wire       [7:0]    dSP_138_b;
  wire       [7:0]    dSP_139_a;
  wire       [7:0]    dSP_139_d;
  wire       [7:0]    dSP_139_b;
  wire       [7:0]    dSP_140_a;
  wire       [7:0]    dSP_140_d;
  wire       [7:0]    dSP_140_b;
  wire       [7:0]    dSP_141_a;
  wire       [7:0]    dSP_141_d;
  wire       [7:0]    dSP_141_b;
  wire       [7:0]    dSP_142_a;
  wire       [7:0]    dSP_142_d;
  wire       [7:0]    dSP_142_b;
  wire       [7:0]    dSP_143_a;
  wire       [7:0]    dSP_143_d;
  wire       [7:0]    dSP_143_b;
  wire       [7:0]    dSP_144_a;
  wire       [7:0]    dSP_144_d;
  wire       [7:0]    dSP_144_b;
  wire       [7:0]    dSP_145_a;
  wire       [7:0]    dSP_145_d;
  wire       [7:0]    dSP_145_b;
  wire       [7:0]    dSP_146_a;
  wire       [7:0]    dSP_146_d;
  wire       [7:0]    dSP_146_b;
  wire       [7:0]    dSP_147_a;
  wire       [7:0]    dSP_147_d;
  wire       [7:0]    dSP_147_b;
  wire       [7:0]    dSP_148_a;
  wire       [7:0]    dSP_148_d;
  wire       [7:0]    dSP_148_b;
  wire       [7:0]    dSP_149_a;
  wire       [7:0]    dSP_149_d;
  wire       [7:0]    dSP_149_b;
  wire       [7:0]    dSP_150_a;
  wire       [7:0]    dSP_150_d;
  wire       [7:0]    dSP_150_b;
  wire       [7:0]    dSP_151_a;
  wire       [7:0]    dSP_151_d;
  wire       [7:0]    dSP_151_b;
  wire       [7:0]    dSP_152_a;
  wire       [7:0]    dSP_152_d;
  wire       [7:0]    dSP_152_b;
  wire       [7:0]    dSP_153_a;
  wire       [7:0]    dSP_153_d;
  wire       [7:0]    dSP_153_b;
  wire       [7:0]    dSP_154_a;
  wire       [7:0]    dSP_154_d;
  wire       [7:0]    dSP_154_b;
  wire       [7:0]    dSP_155_a;
  wire       [7:0]    dSP_155_d;
  wire       [7:0]    dSP_155_b;
  wire       [7:0]    dSP_156_a;
  wire       [7:0]    dSP_156_d;
  wire       [7:0]    dSP_156_b;
  wire       [7:0]    dSP_157_a;
  wire       [7:0]    dSP_157_d;
  wire       [7:0]    dSP_157_b;
  wire       [7:0]    dSP_158_a;
  wire       [7:0]    dSP_158_d;
  wire       [7:0]    dSP_158_b;
  wire       [7:0]    dSP_159_a;
  wire       [7:0]    dSP_159_d;
  wire       [7:0]    dSP_159_b;
  wire       [7:0]    dSP_160_a;
  wire       [7:0]    dSP_160_d;
  wire       [7:0]    dSP_160_b;
  wire       [7:0]    dSP_161_a;
  wire       [7:0]    dSP_161_d;
  wire       [7:0]    dSP_161_b;
  wire       [7:0]    dSP_162_a;
  wire       [7:0]    dSP_162_d;
  wire       [7:0]    dSP_162_b;
  wire       [7:0]    dSP_163_a;
  wire       [7:0]    dSP_163_d;
  wire       [7:0]    dSP_163_b;
  wire       [7:0]    dSP_164_a;
  wire       [7:0]    dSP_164_d;
  wire       [7:0]    dSP_164_b;
  wire       [7:0]    dSP_165_a;
  wire       [7:0]    dSP_165_d;
  wire       [7:0]    dSP_165_b;
  wire       [7:0]    dSP_166_a;
  wire       [7:0]    dSP_166_d;
  wire       [7:0]    dSP_166_b;
  wire       [7:0]    dSP_167_a;
  wire       [7:0]    dSP_167_d;
  wire       [7:0]    dSP_167_b;
  wire       [7:0]    dSP_168_a;
  wire       [7:0]    dSP_168_d;
  wire       [7:0]    dSP_168_b;
  wire       [7:0]    dSP_169_a;
  wire       [7:0]    dSP_169_d;
  wire       [7:0]    dSP_169_b;
  wire       [7:0]    dSP_170_a;
  wire       [7:0]    dSP_170_d;
  wire       [7:0]    dSP_170_b;
  wire       [7:0]    dSP_171_a;
  wire       [7:0]    dSP_171_d;
  wire       [7:0]    dSP_171_b;
  wire       [7:0]    dSP_172_a;
  wire       [7:0]    dSP_172_d;
  wire       [7:0]    dSP_172_b;
  wire       [7:0]    dSP_173_a;
  wire       [7:0]    dSP_173_d;
  wire       [7:0]    dSP_173_b;
  wire       [7:0]    dSP_174_a;
  wire       [7:0]    dSP_174_d;
  wire       [7:0]    dSP_174_b;
  wire       [7:0]    dSP_175_a;
  wire       [7:0]    dSP_175_d;
  wire       [7:0]    dSP_175_b;
  wire       [7:0]    dSP_176_a;
  wire       [7:0]    dSP_176_d;
  wire       [7:0]    dSP_176_b;
  wire       [7:0]    dSP_177_a;
  wire       [7:0]    dSP_177_d;
  wire       [7:0]    dSP_177_b;
  wire       [7:0]    dSP_178_a;
  wire       [7:0]    dSP_178_d;
  wire       [7:0]    dSP_178_b;
  wire       [7:0]    dSP_179_a;
  wire       [7:0]    dSP_179_d;
  wire       [7:0]    dSP_179_b;
  wire       [7:0]    dSP_180_a;
  wire       [7:0]    dSP_180_d;
  wire       [7:0]    dSP_180_b;
  wire       [7:0]    dSP_181_a;
  wire       [7:0]    dSP_181_d;
  wire       [7:0]    dSP_181_b;
  wire       [7:0]    dSP_182_a;
  wire       [7:0]    dSP_182_d;
  wire       [7:0]    dSP_182_b;
  wire       [7:0]    dSP_183_a;
  wire       [7:0]    dSP_183_d;
  wire       [7:0]    dSP_183_b;
  wire       [7:0]    dSP_184_a;
  wire       [7:0]    dSP_184_d;
  wire       [7:0]    dSP_184_b;
  wire       [7:0]    dSP_185_a;
  wire       [7:0]    dSP_185_d;
  wire       [7:0]    dSP_185_b;
  wire       [7:0]    dSP_186_a;
  wire       [7:0]    dSP_186_d;
  wire       [7:0]    dSP_186_b;
  wire       [7:0]    dSP_187_a;
  wire       [7:0]    dSP_187_d;
  wire       [7:0]    dSP_187_b;
  wire       [7:0]    dSP_188_a;
  wire       [7:0]    dSP_188_d;
  wire       [7:0]    dSP_188_b;
  wire       [7:0]    dSP_189_a;
  wire       [7:0]    dSP_189_d;
  wire       [7:0]    dSP_189_b;
  wire       [7:0]    dSP_190_a;
  wire       [7:0]    dSP_190_d;
  wire       [7:0]    dSP_190_b;
  wire       [7:0]    dSP_191_a;
  wire       [7:0]    dSP_191_d;
  wire       [7:0]    dSP_191_b;
  wire       [7:0]    dSP_192_a;
  wire       [7:0]    dSP_192_d;
  wire       [7:0]    dSP_192_b;
  wire       [7:0]    dSP_193_a;
  wire       [7:0]    dSP_193_d;
  wire       [7:0]    dSP_193_b;
  wire       [7:0]    dSP_194_a;
  wire       [7:0]    dSP_194_d;
  wire       [7:0]    dSP_194_b;
  wire       [7:0]    dSP_195_a;
  wire       [7:0]    dSP_195_d;
  wire       [7:0]    dSP_195_b;
  wire       [7:0]    dSP_196_a;
  wire       [7:0]    dSP_196_d;
  wire       [7:0]    dSP_196_b;
  wire       [7:0]    dSP_197_a;
  wire       [7:0]    dSP_197_d;
  wire       [7:0]    dSP_197_b;
  wire       [7:0]    dSP_198_a;
  wire       [7:0]    dSP_198_d;
  wire       [7:0]    dSP_198_b;
  wire       [7:0]    dSP_199_a;
  wire       [7:0]    dSP_199_d;
  wire       [7:0]    dSP_199_b;
  wire       [7:0]    dSP_200_a;
  wire       [7:0]    dSP_200_d;
  wire       [7:0]    dSP_200_b;
  wire       [7:0]    dSP_201_a;
  wire       [7:0]    dSP_201_d;
  wire       [7:0]    dSP_201_b;
  wire       [7:0]    dSP_202_a;
  wire       [7:0]    dSP_202_d;
  wire       [7:0]    dSP_202_b;
  wire       [7:0]    dSP_203_a;
  wire       [7:0]    dSP_203_d;
  wire       [7:0]    dSP_203_b;
  wire       [7:0]    dSP_204_a;
  wire       [7:0]    dSP_204_d;
  wire       [7:0]    dSP_204_b;
  wire       [7:0]    dSP_205_a;
  wire       [7:0]    dSP_205_d;
  wire       [7:0]    dSP_205_b;
  wire       [7:0]    dSP_206_a;
  wire       [7:0]    dSP_206_d;
  wire       [7:0]    dSP_206_b;
  wire       [7:0]    dSP_207_a;
  wire       [7:0]    dSP_207_d;
  wire       [7:0]    dSP_207_b;
  wire       [7:0]    dSP_208_a;
  wire       [7:0]    dSP_208_d;
  wire       [7:0]    dSP_208_b;
  wire       [7:0]    dSP_209_a;
  wire       [7:0]    dSP_209_d;
  wire       [7:0]    dSP_209_b;
  wire       [7:0]    dSP_210_a;
  wire       [7:0]    dSP_210_d;
  wire       [7:0]    dSP_210_b;
  wire       [7:0]    dSP_211_a;
  wire       [7:0]    dSP_211_d;
  wire       [7:0]    dSP_211_b;
  wire       [7:0]    dSP_212_a;
  wire       [7:0]    dSP_212_d;
  wire       [7:0]    dSP_212_b;
  wire       [7:0]    dSP_213_a;
  wire       [7:0]    dSP_213_d;
  wire       [7:0]    dSP_213_b;
  wire       [7:0]    dSP_214_a;
  wire       [7:0]    dSP_214_d;
  wire       [7:0]    dSP_214_b;
  wire       [7:0]    dSP_215_a;
  wire       [7:0]    dSP_215_d;
  wire       [7:0]    dSP_215_b;
  wire       [7:0]    dSP_216_a;
  wire       [7:0]    dSP_216_d;
  wire       [7:0]    dSP_216_b;
  wire       [7:0]    dSP_217_a;
  wire       [7:0]    dSP_217_d;
  wire       [7:0]    dSP_217_b;
  wire       [7:0]    dSP_218_a;
  wire       [7:0]    dSP_218_d;
  wire       [7:0]    dSP_218_b;
  wire       [7:0]    dSP_219_a;
  wire       [7:0]    dSP_219_d;
  wire       [7:0]    dSP_219_b;
  wire       [7:0]    dSP_220_a;
  wire       [7:0]    dSP_220_d;
  wire       [7:0]    dSP_220_b;
  wire       [7:0]    dSP_221_a;
  wire       [7:0]    dSP_221_d;
  wire       [7:0]    dSP_221_b;
  wire       [7:0]    dSP_222_a;
  wire       [7:0]    dSP_222_d;
  wire       [7:0]    dSP_222_b;
  wire       [7:0]    dSP_223_a;
  wire       [7:0]    dSP_223_d;
  wire       [7:0]    dSP_223_b;
  wire       [7:0]    dSP_224_a;
  wire       [7:0]    dSP_224_d;
  wire       [7:0]    dSP_224_b;
  wire       [7:0]    dSP_225_a;
  wire       [7:0]    dSP_225_d;
  wire       [7:0]    dSP_225_b;
  wire       [7:0]    dSP_226_a;
  wire       [7:0]    dSP_226_d;
  wire       [7:0]    dSP_226_b;
  wire       [7:0]    dSP_227_a;
  wire       [7:0]    dSP_227_d;
  wire       [7:0]    dSP_227_b;
  wire       [7:0]    dSP_228_a;
  wire       [7:0]    dSP_228_d;
  wire       [7:0]    dSP_228_b;
  wire       [7:0]    dSP_229_a;
  wire       [7:0]    dSP_229_d;
  wire       [7:0]    dSP_229_b;
  wire       [7:0]    dSP_230_a;
  wire       [7:0]    dSP_230_d;
  wire       [7:0]    dSP_230_b;
  wire       [7:0]    dSP_231_a;
  wire       [7:0]    dSP_231_d;
  wire       [7:0]    dSP_231_b;
  wire       [7:0]    dSP_232_a;
  wire       [7:0]    dSP_232_d;
  wire       [7:0]    dSP_232_b;
  wire       [7:0]    dSP_233_a;
  wire       [7:0]    dSP_233_d;
  wire       [7:0]    dSP_233_b;
  wire       [7:0]    dSP_234_a;
  wire       [7:0]    dSP_234_d;
  wire       [7:0]    dSP_234_b;
  wire       [7:0]    dSP_235_a;
  wire       [7:0]    dSP_235_d;
  wire       [7:0]    dSP_235_b;
  wire       [7:0]    dSP_236_a;
  wire       [7:0]    dSP_236_d;
  wire       [7:0]    dSP_236_b;
  wire       [7:0]    dSP_237_a;
  wire       [7:0]    dSP_237_d;
  wire       [7:0]    dSP_237_b;
  wire       [7:0]    dSP_238_a;
  wire       [7:0]    dSP_238_d;
  wire       [7:0]    dSP_238_b;
  wire       [7:0]    dSP_239_a;
  wire       [7:0]    dSP_239_d;
  wire       [7:0]    dSP_239_b;
  wire       [7:0]    dSP_240_a;
  wire       [7:0]    dSP_240_d;
  wire       [7:0]    dSP_240_b;
  wire       [7:0]    dSP_241_a;
  wire       [7:0]    dSP_241_d;
  wire       [7:0]    dSP_241_b;
  wire       [7:0]    dSP_242_a;
  wire       [7:0]    dSP_242_d;
  wire       [7:0]    dSP_242_b;
  wire       [7:0]    dSP_243_a;
  wire       [7:0]    dSP_243_d;
  wire       [7:0]    dSP_243_b;
  wire       [7:0]    dSP_244_a;
  wire       [7:0]    dSP_244_d;
  wire       [7:0]    dSP_244_b;
  wire       [7:0]    dSP_245_a;
  wire       [7:0]    dSP_245_d;
  wire       [7:0]    dSP_245_b;
  wire       [7:0]    dSP_246_a;
  wire       [7:0]    dSP_246_d;
  wire       [7:0]    dSP_246_b;
  wire       [7:0]    dSP_247_a;
  wire       [7:0]    dSP_247_d;
  wire       [7:0]    dSP_247_b;
  wire       [7:0]    dSP_248_a;
  wire       [7:0]    dSP_248_d;
  wire       [7:0]    dSP_248_b;
  wire       [7:0]    dSP_249_a;
  wire       [7:0]    dSP_249_d;
  wire       [7:0]    dSP_249_b;
  wire       [7:0]    dSP_250_a;
  wire       [7:0]    dSP_250_d;
  wire       [7:0]    dSP_250_b;
  wire       [7:0]    dSP_251_a;
  wire       [7:0]    dSP_251_d;
  wire       [7:0]    dSP_251_b;
  wire       [7:0]    dSP_252_a;
  wire       [7:0]    dSP_252_d;
  wire       [7:0]    dSP_252_b;
  wire       [7:0]    dSP_253_a;
  wire       [7:0]    dSP_253_d;
  wire       [7:0]    dSP_253_b;
  wire       [7:0]    dSP_254_a;
  wire       [7:0]    dSP_254_d;
  wire       [7:0]    dSP_254_b;
  wire       [7:0]    dSP_255_a;
  wire       [7:0]    dSP_255_d;
  wire       [7:0]    dSP_255_b;
  wire       [7:0]    dSP_256_a;
  wire       [7:0]    dSP_256_d;
  wire       [7:0]    dSP_256_b;
  wire       [7:0]    dSP_257_a;
  wire       [7:0]    dSP_257_d;
  wire       [7:0]    dSP_257_b;
  wire       [7:0]    dSP_258_a;
  wire       [7:0]    dSP_258_d;
  wire       [7:0]    dSP_258_b;
  wire       [7:0]    dSP_259_a;
  wire       [7:0]    dSP_259_d;
  wire       [7:0]    dSP_259_b;
  wire       [7:0]    dSP_260_a;
  wire       [7:0]    dSP_260_d;
  wire       [7:0]    dSP_260_b;
  wire       [7:0]    dSP_261_a;
  wire       [7:0]    dSP_261_d;
  wire       [7:0]    dSP_261_b;
  wire       [7:0]    dSP_262_a;
  wire       [7:0]    dSP_262_d;
  wire       [7:0]    dSP_262_b;
  wire       [7:0]    dSP_263_a;
  wire       [7:0]    dSP_263_d;
  wire       [7:0]    dSP_263_b;
  wire       [7:0]    dSP_264_a;
  wire       [7:0]    dSP_264_d;
  wire       [7:0]    dSP_264_b;
  wire       [7:0]    dSP_265_a;
  wire       [7:0]    dSP_265_d;
  wire       [7:0]    dSP_265_b;
  wire       [7:0]    dSP_266_a;
  wire       [7:0]    dSP_266_d;
  wire       [7:0]    dSP_266_b;
  wire       [7:0]    dSP_267_a;
  wire       [7:0]    dSP_267_d;
  wire       [7:0]    dSP_267_b;
  wire       [7:0]    dSP_268_a;
  wire       [7:0]    dSP_268_d;
  wire       [7:0]    dSP_268_b;
  wire       [7:0]    dSP_269_a;
  wire       [7:0]    dSP_269_d;
  wire       [7:0]    dSP_269_b;
  wire       [7:0]    dSP_270_a;
  wire       [7:0]    dSP_270_d;
  wire       [7:0]    dSP_270_b;
  wire       [7:0]    dSP_271_a;
  wire       [7:0]    dSP_271_d;
  wire       [7:0]    dSP_271_b;
  wire       [7:0]    dSP_272_a;
  wire       [7:0]    dSP_272_d;
  wire       [7:0]    dSP_272_b;
  wire       [7:0]    dSP_273_a;
  wire       [7:0]    dSP_273_d;
  wire       [7:0]    dSP_273_b;
  wire       [7:0]    dSP_274_a;
  wire       [7:0]    dSP_274_d;
  wire       [7:0]    dSP_274_b;
  wire       [7:0]    dSP_275_a;
  wire       [7:0]    dSP_275_d;
  wire       [7:0]    dSP_275_b;
  wire       [7:0]    dSP_276_a;
  wire       [7:0]    dSP_276_d;
  wire       [7:0]    dSP_276_b;
  wire       [7:0]    dSP_277_a;
  wire       [7:0]    dSP_277_d;
  wire       [7:0]    dSP_277_b;
  wire       [7:0]    dSP_278_a;
  wire       [7:0]    dSP_278_d;
  wire       [7:0]    dSP_278_b;
  wire       [7:0]    dSP_279_a;
  wire       [7:0]    dSP_279_d;
  wire       [7:0]    dSP_279_b;
  wire       [7:0]    dSP_280_a;
  wire       [7:0]    dSP_280_d;
  wire       [7:0]    dSP_280_b;
  wire       [7:0]    dSP_281_a;
  wire       [7:0]    dSP_281_d;
  wire       [7:0]    dSP_281_b;
  wire       [7:0]    dSP_282_a;
  wire       [7:0]    dSP_282_d;
  wire       [7:0]    dSP_282_b;
  wire       [7:0]    dSP_283_a;
  wire       [7:0]    dSP_283_d;
  wire       [7:0]    dSP_283_b;
  wire       [7:0]    dSP_284_a;
  wire       [7:0]    dSP_284_d;
  wire       [7:0]    dSP_284_b;
  wire       [7:0]    dSP_285_a;
  wire       [7:0]    dSP_285_d;
  wire       [7:0]    dSP_285_b;
  wire       [7:0]    dSP_286_a;
  wire       [7:0]    dSP_286_d;
  wire       [7:0]    dSP_286_b;
  wire       [7:0]    dSP_287_a;
  wire       [7:0]    dSP_287_d;
  wire       [7:0]    dSP_287_b;
  wire       [7:0]    dSP_288_a;
  wire       [7:0]    dSP_288_d;
  wire       [7:0]    dSP_288_b;
  wire       [7:0]    dSP_289_a;
  wire       [7:0]    dSP_289_d;
  wire       [7:0]    dSP_289_b;
  wire       [7:0]    dSP_290_a;
  wire       [7:0]    dSP_290_d;
  wire       [7:0]    dSP_290_b;
  wire       [7:0]    dSP_291_a;
  wire       [7:0]    dSP_291_d;
  wire       [7:0]    dSP_291_b;
  wire       [7:0]    dSP_292_a;
  wire       [7:0]    dSP_292_d;
  wire       [7:0]    dSP_292_b;
  wire       [7:0]    dSP_293_a;
  wire       [7:0]    dSP_293_d;
  wire       [7:0]    dSP_293_b;
  wire       [7:0]    dSP_294_a;
  wire       [7:0]    dSP_294_d;
  wire       [7:0]    dSP_294_b;
  wire       [7:0]    dSP_295_a;
  wire       [7:0]    dSP_295_d;
  wire       [7:0]    dSP_295_b;
  wire       [7:0]    dSP_296_a;
  wire       [7:0]    dSP_296_d;
  wire       [7:0]    dSP_296_b;
  wire       [7:0]    dSP_297_a;
  wire       [7:0]    dSP_297_d;
  wire       [7:0]    dSP_297_b;
  wire       [7:0]    dSP_298_a;
  wire       [7:0]    dSP_298_d;
  wire       [7:0]    dSP_298_b;
  wire       [7:0]    dSP_299_a;
  wire       [7:0]    dSP_299_d;
  wire       [7:0]    dSP_299_b;
  wire       [7:0]    dSP_300_a;
  wire       [7:0]    dSP_300_d;
  wire       [7:0]    dSP_300_b;
  wire       [7:0]    dSP_301_a;
  wire       [7:0]    dSP_301_d;
  wire       [7:0]    dSP_301_b;
  wire       [7:0]    dSP_302_a;
  wire       [7:0]    dSP_302_d;
  wire       [7:0]    dSP_302_b;
  wire       [7:0]    dSP_303_a;
  wire       [7:0]    dSP_303_d;
  wire       [7:0]    dSP_303_b;
  wire       [7:0]    dSP_304_a;
  wire       [7:0]    dSP_304_d;
  wire       [7:0]    dSP_304_b;
  wire       [7:0]    dSP_305_a;
  wire       [7:0]    dSP_305_d;
  wire       [7:0]    dSP_305_b;
  wire       [7:0]    dSP_306_a;
  wire       [7:0]    dSP_306_d;
  wire       [7:0]    dSP_306_b;
  wire       [7:0]    dSP_307_a;
  wire       [7:0]    dSP_307_d;
  wire       [7:0]    dSP_307_b;
  wire       [7:0]    dSP_308_a;
  wire       [7:0]    dSP_308_d;
  wire       [7:0]    dSP_308_b;
  wire       [7:0]    dSP_309_a;
  wire       [7:0]    dSP_309_d;
  wire       [7:0]    dSP_309_b;
  wire       [7:0]    dSP_310_a;
  wire       [7:0]    dSP_310_d;
  wire       [7:0]    dSP_310_b;
  wire       [7:0]    dSP_311_a;
  wire       [7:0]    dSP_311_d;
  wire       [7:0]    dSP_311_b;
  wire       [7:0]    dSP_312_a;
  wire       [7:0]    dSP_312_d;
  wire       [7:0]    dSP_312_b;
  wire       [7:0]    dSP_313_a;
  wire       [7:0]    dSP_313_d;
  wire       [7:0]    dSP_313_b;
  wire       [7:0]    dSP_314_a;
  wire       [7:0]    dSP_314_d;
  wire       [7:0]    dSP_314_b;
  wire       [7:0]    dSP_315_a;
  wire       [7:0]    dSP_315_d;
  wire       [7:0]    dSP_315_b;
  wire       [7:0]    dSP_316_a;
  wire       [7:0]    dSP_316_d;
  wire       [7:0]    dSP_316_b;
  wire       [7:0]    dSP_317_a;
  wire       [7:0]    dSP_317_d;
  wire       [7:0]    dSP_317_b;
  wire       [7:0]    dSP_318_a;
  wire       [7:0]    dSP_318_d;
  wire       [7:0]    dSP_318_b;
  wire       [7:0]    dSP_319_a;
  wire       [7:0]    dSP_319_d;
  wire       [7:0]    dSP_319_b;
  wire       [7:0]    dSP_320_a;
  wire       [7:0]    dSP_320_d;
  wire       [7:0]    dSP_320_b;
  wire       [7:0]    dSP_321_a;
  wire       [7:0]    dSP_321_d;
  wire       [7:0]    dSP_321_b;
  wire       [7:0]    dSP_322_a;
  wire       [7:0]    dSP_322_d;
  wire       [7:0]    dSP_322_b;
  wire       [7:0]    dSP_323_a;
  wire       [7:0]    dSP_323_d;
  wire       [7:0]    dSP_323_b;
  wire       [7:0]    dSP_324_a;
  wire       [7:0]    dSP_324_d;
  wire       [7:0]    dSP_324_b;
  wire       [7:0]    dSP_325_a;
  wire       [7:0]    dSP_325_d;
  wire       [7:0]    dSP_325_b;
  wire       [7:0]    dSP_326_a;
  wire       [7:0]    dSP_326_d;
  wire       [7:0]    dSP_326_b;
  wire       [7:0]    dSP_327_a;
  wire       [7:0]    dSP_327_d;
  wire       [7:0]    dSP_327_b;
  wire       [7:0]    dSP_328_a;
  wire       [7:0]    dSP_328_d;
  wire       [7:0]    dSP_328_b;
  wire       [7:0]    dSP_329_a;
  wire       [7:0]    dSP_329_d;
  wire       [7:0]    dSP_329_b;
  wire       [7:0]    dSP_330_a;
  wire       [7:0]    dSP_330_d;
  wire       [7:0]    dSP_330_b;
  wire       [7:0]    dSP_331_a;
  wire       [7:0]    dSP_331_d;
  wire       [7:0]    dSP_331_b;
  wire       [7:0]    dSP_332_a;
  wire       [7:0]    dSP_332_d;
  wire       [7:0]    dSP_332_b;
  wire       [7:0]    dSP_333_a;
  wire       [7:0]    dSP_333_d;
  wire       [7:0]    dSP_333_b;
  wire       [7:0]    dSP_334_a;
  wire       [7:0]    dSP_334_d;
  wire       [7:0]    dSP_334_b;
  wire       [7:0]    dSP_335_a;
  wire       [7:0]    dSP_335_d;
  wire       [7:0]    dSP_335_b;
  wire       [7:0]    dSP_336_a;
  wire       [7:0]    dSP_336_d;
  wire       [7:0]    dSP_336_b;
  wire       [7:0]    dSP_337_a;
  wire       [7:0]    dSP_337_d;
  wire       [7:0]    dSP_337_b;
  wire       [7:0]    dSP_338_a;
  wire       [7:0]    dSP_338_d;
  wire       [7:0]    dSP_338_b;
  wire       [7:0]    dSP_339_a;
  wire       [7:0]    dSP_339_d;
  wire       [7:0]    dSP_339_b;
  wire       [7:0]    dSP_340_a;
  wire       [7:0]    dSP_340_d;
  wire       [7:0]    dSP_340_b;
  wire       [7:0]    dSP_341_a;
  wire       [7:0]    dSP_341_d;
  wire       [7:0]    dSP_341_b;
  wire       [7:0]    dSP_342_a;
  wire       [7:0]    dSP_342_d;
  wire       [7:0]    dSP_342_b;
  wire       [7:0]    dSP_343_a;
  wire       [7:0]    dSP_343_d;
  wire       [7:0]    dSP_343_b;
  wire       [7:0]    dSP_344_a;
  wire       [7:0]    dSP_344_d;
  wire       [7:0]    dSP_344_b;
  wire       [7:0]    dSP_345_a;
  wire       [7:0]    dSP_345_d;
  wire       [7:0]    dSP_345_b;
  wire       [7:0]    dSP_346_a;
  wire       [7:0]    dSP_346_d;
  wire       [7:0]    dSP_346_b;
  wire       [7:0]    dSP_347_a;
  wire       [7:0]    dSP_347_d;
  wire       [7:0]    dSP_347_b;
  wire       [7:0]    dSP_348_a;
  wire       [7:0]    dSP_348_d;
  wire       [7:0]    dSP_348_b;
  wire       [7:0]    dSP_349_a;
  wire       [7:0]    dSP_349_d;
  wire       [7:0]    dSP_349_b;
  wire       [7:0]    dSP_350_a;
  wire       [7:0]    dSP_350_d;
  wire       [7:0]    dSP_350_b;
  wire       [7:0]    dSP_351_a;
  wire       [7:0]    dSP_351_d;
  wire       [7:0]    dSP_351_b;
  wire       [7:0]    dSP_352_a;
  wire       [7:0]    dSP_352_d;
  wire       [7:0]    dSP_352_b;
  wire       [7:0]    dSP_353_a;
  wire       [7:0]    dSP_353_d;
  wire       [7:0]    dSP_353_b;
  wire       [7:0]    dSP_354_a;
  wire       [7:0]    dSP_354_d;
  wire       [7:0]    dSP_354_b;
  wire       [7:0]    dSP_355_a;
  wire       [7:0]    dSP_355_d;
  wire       [7:0]    dSP_355_b;
  wire       [7:0]    dSP_356_a;
  wire       [7:0]    dSP_356_d;
  wire       [7:0]    dSP_356_b;
  wire       [7:0]    dSP_357_a;
  wire       [7:0]    dSP_357_d;
  wire       [7:0]    dSP_357_b;
  wire       [7:0]    dSP_358_a;
  wire       [7:0]    dSP_358_d;
  wire       [7:0]    dSP_358_b;
  wire       [7:0]    dSP_359_a;
  wire       [7:0]    dSP_359_d;
  wire       [7:0]    dSP_359_b;
  wire       [7:0]    dSP_360_a;
  wire       [7:0]    dSP_360_d;
  wire       [7:0]    dSP_360_b;
  wire       [7:0]    dSP_361_a;
  wire       [7:0]    dSP_361_d;
  wire       [7:0]    dSP_361_b;
  wire       [7:0]    dSP_362_a;
  wire       [7:0]    dSP_362_d;
  wire       [7:0]    dSP_362_b;
  wire       [7:0]    dSP_363_a;
  wire       [7:0]    dSP_363_d;
  wire       [7:0]    dSP_363_b;
  wire       [7:0]    dSP_364_a;
  wire       [7:0]    dSP_364_d;
  wire       [7:0]    dSP_364_b;
  wire       [7:0]    dSP_365_a;
  wire       [7:0]    dSP_365_d;
  wire       [7:0]    dSP_365_b;
  wire       [7:0]    dSP_366_a;
  wire       [7:0]    dSP_366_d;
  wire       [7:0]    dSP_366_b;
  wire       [7:0]    dSP_367_a;
  wire       [7:0]    dSP_367_d;
  wire       [7:0]    dSP_367_b;
  wire       [7:0]    dSP_368_a;
  wire       [7:0]    dSP_368_d;
  wire       [7:0]    dSP_368_b;
  wire       [7:0]    dSP_369_a;
  wire       [7:0]    dSP_369_d;
  wire       [7:0]    dSP_369_b;
  wire       [7:0]    dSP_370_a;
  wire       [7:0]    dSP_370_d;
  wire       [7:0]    dSP_370_b;
  wire       [7:0]    dSP_371_a;
  wire       [7:0]    dSP_371_d;
  wire       [7:0]    dSP_371_b;
  wire       [7:0]    dSP_372_a;
  wire       [7:0]    dSP_372_d;
  wire       [7:0]    dSP_372_b;
  wire       [7:0]    dSP_373_a;
  wire       [7:0]    dSP_373_d;
  wire       [7:0]    dSP_373_b;
  wire       [7:0]    dSP_374_a;
  wire       [7:0]    dSP_374_d;
  wire       [7:0]    dSP_374_b;
  wire       [7:0]    dSP_375_a;
  wire       [7:0]    dSP_375_d;
  wire       [7:0]    dSP_375_b;
  wire       [7:0]    dSP_376_a;
  wire       [7:0]    dSP_376_d;
  wire       [7:0]    dSP_376_b;
  wire       [7:0]    dSP_377_a;
  wire       [7:0]    dSP_377_d;
  wire       [7:0]    dSP_377_b;
  wire       [7:0]    dSP_378_a;
  wire       [7:0]    dSP_378_d;
  wire       [7:0]    dSP_378_b;
  wire       [7:0]    dSP_379_a;
  wire       [7:0]    dSP_379_d;
  wire       [7:0]    dSP_379_b;
  wire       [7:0]    dSP_380_a;
  wire       [7:0]    dSP_380_d;
  wire       [7:0]    dSP_380_b;
  wire       [7:0]    dSP_381_a;
  wire       [7:0]    dSP_381_d;
  wire       [7:0]    dSP_381_b;
  wire       [7:0]    dSP_382_a;
  wire       [7:0]    dSP_382_d;
  wire       [7:0]    dSP_382_b;
  wire       [7:0]    dSP_383_a;
  wire       [7:0]    dSP_383_d;
  wire       [7:0]    dSP_383_b;
  wire       [7:0]    dSP_384_a;
  wire       [7:0]    dSP_384_d;
  wire       [7:0]    dSP_384_b;
  wire       [7:0]    dSP_385_a;
  wire       [7:0]    dSP_385_d;
  wire       [7:0]    dSP_385_b;
  wire       [7:0]    dSP_386_a;
  wire       [7:0]    dSP_386_d;
  wire       [7:0]    dSP_386_b;
  wire       [7:0]    dSP_387_a;
  wire       [7:0]    dSP_387_d;
  wire       [7:0]    dSP_387_b;
  wire       [7:0]    dSP_388_a;
  wire       [7:0]    dSP_388_d;
  wire       [7:0]    dSP_388_b;
  wire       [7:0]    dSP_389_a;
  wire       [7:0]    dSP_389_d;
  wire       [7:0]    dSP_389_b;
  wire       [7:0]    dSP_390_a;
  wire       [7:0]    dSP_390_d;
  wire       [7:0]    dSP_390_b;
  wire       [7:0]    dSP_391_a;
  wire       [7:0]    dSP_391_d;
  wire       [7:0]    dSP_391_b;
  wire       [7:0]    dSP_392_a;
  wire       [7:0]    dSP_392_d;
  wire       [7:0]    dSP_392_b;
  wire       [7:0]    dSP_393_a;
  wire       [7:0]    dSP_393_d;
  wire       [7:0]    dSP_393_b;
  wire       [7:0]    dSP_394_a;
  wire       [7:0]    dSP_394_d;
  wire       [7:0]    dSP_394_b;
  wire       [7:0]    dSP_395_a;
  wire       [7:0]    dSP_395_d;
  wire       [7:0]    dSP_395_b;
  wire       [7:0]    dSP_396_a;
  wire       [7:0]    dSP_396_d;
  wire       [7:0]    dSP_396_b;
  wire       [7:0]    dSP_397_a;
  wire       [7:0]    dSP_397_d;
  wire       [7:0]    dSP_397_b;
  wire       [7:0]    dSP_398_a;
  wire       [7:0]    dSP_398_d;
  wire       [7:0]    dSP_398_b;
  wire       [7:0]    dSP_399_a;
  wire       [7:0]    dSP_399_d;
  wire       [7:0]    dSP_399_b;
  wire       [7:0]    dSP_400_a;
  wire       [7:0]    dSP_400_d;
  wire       [7:0]    dSP_400_b;
  wire       [7:0]    dSP_401_a;
  wire       [7:0]    dSP_401_d;
  wire       [7:0]    dSP_401_b;
  wire       [7:0]    dSP_402_a;
  wire       [7:0]    dSP_402_d;
  wire       [7:0]    dSP_402_b;
  wire       [7:0]    dSP_403_a;
  wire       [7:0]    dSP_403_d;
  wire       [7:0]    dSP_403_b;
  wire       [7:0]    dSP_404_a;
  wire       [7:0]    dSP_404_d;
  wire       [7:0]    dSP_404_b;
  wire       [7:0]    dSP_405_a;
  wire       [7:0]    dSP_405_d;
  wire       [7:0]    dSP_405_b;
  wire       [7:0]    dSP_406_a;
  wire       [7:0]    dSP_406_d;
  wire       [7:0]    dSP_406_b;
  wire       [7:0]    dSP_407_a;
  wire       [7:0]    dSP_407_d;
  wire       [7:0]    dSP_407_b;
  wire       [7:0]    dSP_408_a;
  wire       [7:0]    dSP_408_d;
  wire       [7:0]    dSP_408_b;
  wire       [7:0]    dSP_409_a;
  wire       [7:0]    dSP_409_d;
  wire       [7:0]    dSP_409_b;
  wire       [7:0]    dSP_410_a;
  wire       [7:0]    dSP_410_d;
  wire       [7:0]    dSP_410_b;
  wire       [7:0]    dSP_411_a;
  wire       [7:0]    dSP_411_d;
  wire       [7:0]    dSP_411_b;
  wire       [7:0]    dSP_412_a;
  wire       [7:0]    dSP_412_d;
  wire       [7:0]    dSP_412_b;
  wire       [7:0]    dSP_413_a;
  wire       [7:0]    dSP_413_d;
  wire       [7:0]    dSP_413_b;
  wire       [7:0]    dSP_414_a;
  wire       [7:0]    dSP_414_d;
  wire       [7:0]    dSP_414_b;
  wire       [7:0]    dSP_415_a;
  wire       [7:0]    dSP_415_d;
  wire       [7:0]    dSP_415_b;
  wire       [7:0]    dSP_416_a;
  wire       [7:0]    dSP_416_d;
  wire       [7:0]    dSP_416_b;
  wire       [7:0]    dSP_417_a;
  wire       [7:0]    dSP_417_d;
  wire       [7:0]    dSP_417_b;
  wire       [7:0]    dSP_418_a;
  wire       [7:0]    dSP_418_d;
  wire       [7:0]    dSP_418_b;
  wire       [7:0]    dSP_419_a;
  wire       [7:0]    dSP_419_d;
  wire       [7:0]    dSP_419_b;
  wire       [7:0]    dSP_420_a;
  wire       [7:0]    dSP_420_d;
  wire       [7:0]    dSP_420_b;
  wire       [7:0]    dSP_421_a;
  wire       [7:0]    dSP_421_d;
  wire       [7:0]    dSP_421_b;
  wire       [7:0]    dSP_422_a;
  wire       [7:0]    dSP_422_d;
  wire       [7:0]    dSP_422_b;
  wire       [7:0]    dSP_423_a;
  wire       [7:0]    dSP_423_d;
  wire       [7:0]    dSP_423_b;
  wire       [7:0]    dSP_424_a;
  wire       [7:0]    dSP_424_d;
  wire       [7:0]    dSP_424_b;
  wire       [7:0]    dSP_425_a;
  wire       [7:0]    dSP_425_d;
  wire       [7:0]    dSP_425_b;
  wire       [7:0]    dSP_426_a;
  wire       [7:0]    dSP_426_d;
  wire       [7:0]    dSP_426_b;
  wire       [7:0]    dSP_427_a;
  wire       [7:0]    dSP_427_d;
  wire       [7:0]    dSP_427_b;
  wire       [7:0]    dSP_428_a;
  wire       [7:0]    dSP_428_d;
  wire       [7:0]    dSP_428_b;
  wire       [7:0]    dSP_429_a;
  wire       [7:0]    dSP_429_d;
  wire       [7:0]    dSP_429_b;
  wire       [7:0]    dSP_430_a;
  wire       [7:0]    dSP_430_d;
  wire       [7:0]    dSP_430_b;
  wire       [7:0]    dSP_431_a;
  wire       [7:0]    dSP_431_d;
  wire       [7:0]    dSP_431_b;
  wire       [7:0]    dSP_432_a;
  wire       [7:0]    dSP_432_d;
  wire       [7:0]    dSP_432_b;
  wire       [7:0]    dSP_433_a;
  wire       [7:0]    dSP_433_d;
  wire       [7:0]    dSP_433_b;
  wire       [7:0]    dSP_434_a;
  wire       [7:0]    dSP_434_d;
  wire       [7:0]    dSP_434_b;
  wire       [7:0]    dSP_435_a;
  wire       [7:0]    dSP_435_d;
  wire       [7:0]    dSP_435_b;
  wire       [7:0]    dSP_436_a;
  wire       [7:0]    dSP_436_d;
  wire       [7:0]    dSP_436_b;
  wire       [7:0]    dSP_437_a;
  wire       [7:0]    dSP_437_d;
  wire       [7:0]    dSP_437_b;
  wire       [7:0]    dSP_438_a;
  wire       [7:0]    dSP_438_d;
  wire       [7:0]    dSP_438_b;
  wire       [7:0]    dSP_439_a;
  wire       [7:0]    dSP_439_d;
  wire       [7:0]    dSP_439_b;
  wire       [7:0]    dSP_440_a;
  wire       [7:0]    dSP_440_d;
  wire       [7:0]    dSP_440_b;
  wire       [7:0]    dSP_441_a;
  wire       [7:0]    dSP_441_d;
  wire       [7:0]    dSP_441_b;
  wire       [7:0]    dSP_442_a;
  wire       [7:0]    dSP_442_d;
  wire       [7:0]    dSP_442_b;
  wire       [7:0]    dSP_443_a;
  wire       [7:0]    dSP_443_d;
  wire       [7:0]    dSP_443_b;
  wire       [7:0]    dSP_444_a;
  wire       [7:0]    dSP_444_d;
  wire       [7:0]    dSP_444_b;
  wire       [7:0]    dSP_445_a;
  wire       [7:0]    dSP_445_d;
  wire       [7:0]    dSP_445_b;
  wire       [7:0]    dSP_446_a;
  wire       [7:0]    dSP_446_d;
  wire       [7:0]    dSP_446_b;
  wire       [7:0]    dSP_447_a;
  wire       [7:0]    dSP_447_d;
  wire       [7:0]    dSP_447_b;
  wire       [7:0]    dSP_448_a;
  wire       [7:0]    dSP_448_d;
  wire       [7:0]    dSP_448_b;
  wire       [7:0]    dSP_449_a;
  wire       [7:0]    dSP_449_d;
  wire       [7:0]    dSP_449_b;
  wire       [7:0]    dSP_450_a;
  wire       [7:0]    dSP_450_d;
  wire       [7:0]    dSP_450_b;
  wire       [7:0]    dSP_451_a;
  wire       [7:0]    dSP_451_d;
  wire       [7:0]    dSP_451_b;
  wire       [7:0]    dSP_452_a;
  wire       [7:0]    dSP_452_d;
  wire       [7:0]    dSP_452_b;
  wire       [7:0]    dSP_453_a;
  wire       [7:0]    dSP_453_d;
  wire       [7:0]    dSP_453_b;
  wire       [7:0]    dSP_454_a;
  wire       [7:0]    dSP_454_d;
  wire       [7:0]    dSP_454_b;
  wire       [7:0]    dSP_455_a;
  wire       [7:0]    dSP_455_d;
  wire       [7:0]    dSP_455_b;
  wire       [7:0]    dSP_456_a;
  wire       [7:0]    dSP_456_d;
  wire       [7:0]    dSP_456_b;
  wire       [7:0]    dSP_457_a;
  wire       [7:0]    dSP_457_d;
  wire       [7:0]    dSP_457_b;
  wire       [7:0]    dSP_458_a;
  wire       [7:0]    dSP_458_d;
  wire       [7:0]    dSP_458_b;
  wire       [7:0]    dSP_459_a;
  wire       [7:0]    dSP_459_d;
  wire       [7:0]    dSP_459_b;
  wire       [7:0]    dSP_460_a;
  wire       [7:0]    dSP_460_d;
  wire       [7:0]    dSP_460_b;
  wire       [7:0]    dSP_461_a;
  wire       [7:0]    dSP_461_d;
  wire       [7:0]    dSP_461_b;
  wire       [7:0]    dSP_462_a;
  wire       [7:0]    dSP_462_d;
  wire       [7:0]    dSP_462_b;
  wire       [7:0]    dSP_463_a;
  wire       [7:0]    dSP_463_d;
  wire       [7:0]    dSP_463_b;
  wire       [7:0]    dSP_464_a;
  wire       [7:0]    dSP_464_d;
  wire       [7:0]    dSP_464_b;
  wire       [7:0]    dSP_465_a;
  wire       [7:0]    dSP_465_d;
  wire       [7:0]    dSP_465_b;
  wire       [7:0]    dSP_466_a;
  wire       [7:0]    dSP_466_d;
  wire       [7:0]    dSP_466_b;
  wire       [7:0]    dSP_467_a;
  wire       [7:0]    dSP_467_d;
  wire       [7:0]    dSP_467_b;
  wire       [7:0]    dSP_468_a;
  wire       [7:0]    dSP_468_d;
  wire       [7:0]    dSP_468_b;
  wire       [7:0]    dSP_469_a;
  wire       [7:0]    dSP_469_d;
  wire       [7:0]    dSP_469_b;
  wire       [7:0]    dSP_470_a;
  wire       [7:0]    dSP_470_d;
  wire       [7:0]    dSP_470_b;
  wire       [7:0]    dSP_471_a;
  wire       [7:0]    dSP_471_d;
  wire       [7:0]    dSP_471_b;
  wire       [7:0]    dSP_472_a;
  wire       [7:0]    dSP_472_d;
  wire       [7:0]    dSP_472_b;
  wire       [7:0]    dSP_473_a;
  wire       [7:0]    dSP_473_d;
  wire       [7:0]    dSP_473_b;
  wire       [7:0]    dSP_474_a;
  wire       [7:0]    dSP_474_d;
  wire       [7:0]    dSP_474_b;
  wire       [7:0]    dSP_475_a;
  wire       [7:0]    dSP_475_d;
  wire       [7:0]    dSP_475_b;
  wire       [7:0]    dSP_476_a;
  wire       [7:0]    dSP_476_d;
  wire       [7:0]    dSP_476_b;
  wire       [7:0]    dSP_477_a;
  wire       [7:0]    dSP_477_d;
  wire       [7:0]    dSP_477_b;
  wire       [7:0]    dSP_478_a;
  wire       [7:0]    dSP_478_d;
  wire       [7:0]    dSP_478_b;
  wire       [7:0]    dSP_479_a;
  wire       [7:0]    dSP_479_d;
  wire       [7:0]    dSP_479_b;
  wire       [7:0]    dSP_480_a;
  wire       [7:0]    dSP_480_d;
  wire       [7:0]    dSP_480_b;
  wire       [7:0]    dSP_481_a;
  wire       [7:0]    dSP_481_d;
  wire       [7:0]    dSP_481_b;
  wire       [7:0]    dSP_482_a;
  wire       [7:0]    dSP_482_d;
  wire       [7:0]    dSP_482_b;
  wire       [7:0]    dSP_483_a;
  wire       [7:0]    dSP_483_d;
  wire       [7:0]    dSP_483_b;
  wire       [7:0]    dSP_484_a;
  wire       [7:0]    dSP_484_d;
  wire       [7:0]    dSP_484_b;
  wire       [7:0]    dSP_485_a;
  wire       [7:0]    dSP_485_d;
  wire       [7:0]    dSP_485_b;
  wire       [7:0]    dSP_486_a;
  wire       [7:0]    dSP_486_d;
  wire       [7:0]    dSP_486_b;
  wire       [7:0]    dSP_487_a;
  wire       [7:0]    dSP_487_d;
  wire       [7:0]    dSP_487_b;
  wire       [7:0]    dSP_488_a;
  wire       [7:0]    dSP_488_d;
  wire       [7:0]    dSP_488_b;
  wire       [7:0]    dSP_489_a;
  wire       [7:0]    dSP_489_d;
  wire       [7:0]    dSP_489_b;
  wire       [7:0]    dSP_490_a;
  wire       [7:0]    dSP_490_d;
  wire       [7:0]    dSP_490_b;
  wire       [7:0]    dSP_491_a;
  wire       [7:0]    dSP_491_d;
  wire       [7:0]    dSP_491_b;
  wire       [7:0]    dSP_492_a;
  wire       [7:0]    dSP_492_d;
  wire       [7:0]    dSP_492_b;
  wire       [7:0]    dSP_493_a;
  wire       [7:0]    dSP_493_d;
  wire       [7:0]    dSP_493_b;
  wire       [7:0]    dSP_494_a;
  wire       [7:0]    dSP_494_d;
  wire       [7:0]    dSP_494_b;
  wire       [7:0]    dSP_495_a;
  wire       [7:0]    dSP_495_d;
  wire       [7:0]    dSP_495_b;
  wire       [7:0]    dSP_496_a;
  wire       [7:0]    dSP_496_d;
  wire       [7:0]    dSP_496_b;
  wire       [7:0]    dSP_497_a;
  wire       [7:0]    dSP_497_d;
  wire       [7:0]    dSP_497_b;
  wire       [7:0]    dSP_498_a;
  wire       [7:0]    dSP_498_d;
  wire       [7:0]    dSP_498_b;
  wire       [7:0]    dSP_499_a;
  wire       [7:0]    dSP_499_d;
  wire       [7:0]    dSP_499_b;
  wire       [7:0]    dSP_500_a;
  wire       [7:0]    dSP_500_d;
  wire       [7:0]    dSP_500_b;
  wire       [7:0]    dSP_501_a;
  wire       [7:0]    dSP_501_d;
  wire       [7:0]    dSP_501_b;
  wire       [7:0]    dSP_502_a;
  wire       [7:0]    dSP_502_d;
  wire       [7:0]    dSP_502_b;
  wire       [7:0]    dSP_503_a;
  wire       [7:0]    dSP_503_d;
  wire       [7:0]    dSP_503_b;
  wire       [7:0]    dSP_504_a;
  wire       [7:0]    dSP_504_d;
  wire       [7:0]    dSP_504_b;
  wire       [7:0]    dSP_505_a;
  wire       [7:0]    dSP_505_d;
  wire       [7:0]    dSP_505_b;
  wire       [7:0]    dSP_506_a;
  wire       [7:0]    dSP_506_d;
  wire       [7:0]    dSP_506_b;
  wire       [7:0]    dSP_507_a;
  wire       [7:0]    dSP_507_d;
  wire       [7:0]    dSP_507_b;
  wire       [7:0]    dSP_508_a;
  wire       [7:0]    dSP_508_d;
  wire       [7:0]    dSP_508_b;
  wire       [7:0]    dSP_509_a;
  wire       [7:0]    dSP_509_d;
  wire       [7:0]    dSP_509_b;
  wire       [7:0]    dSP_510_a;
  wire       [7:0]    dSP_510_d;
  wire       [7:0]    dSP_510_b;
  wire       [7:0]    dSP_511_a;
  wire       [7:0]    dSP_511_d;
  wire       [7:0]    dSP_511_b;
  wire       [7:0]    dSP_512_a;
  wire       [7:0]    dSP_512_d;
  wire       [7:0]    dSP_512_b;
  wire       [7:0]    dSP_513_a;
  wire       [7:0]    dSP_513_d;
  wire       [7:0]    dSP_513_b;
  wire       [7:0]    dSP_514_a;
  wire       [7:0]    dSP_514_d;
  wire       [7:0]    dSP_514_b;
  wire       [7:0]    dSP_515_a;
  wire       [7:0]    dSP_515_d;
  wire       [7:0]    dSP_515_b;
  wire       [7:0]    dSP_516_a;
  wire       [7:0]    dSP_516_d;
  wire       [7:0]    dSP_516_b;
  wire       [7:0]    dSP_517_a;
  wire       [7:0]    dSP_517_d;
  wire       [7:0]    dSP_517_b;
  wire       [7:0]    dSP_518_a;
  wire       [7:0]    dSP_518_d;
  wire       [7:0]    dSP_518_b;
  wire       [7:0]    dSP_519_a;
  wire       [7:0]    dSP_519_d;
  wire       [7:0]    dSP_519_b;
  wire       [7:0]    dSP_520_a;
  wire       [7:0]    dSP_520_d;
  wire       [7:0]    dSP_520_b;
  wire       [7:0]    dSP_521_a;
  wire       [7:0]    dSP_521_d;
  wire       [7:0]    dSP_521_b;
  wire       [7:0]    dSP_522_a;
  wire       [7:0]    dSP_522_d;
  wire       [7:0]    dSP_522_b;
  wire       [7:0]    dSP_523_a;
  wire       [7:0]    dSP_523_d;
  wire       [7:0]    dSP_523_b;
  wire       [7:0]    dSP_524_a;
  wire       [7:0]    dSP_524_d;
  wire       [7:0]    dSP_524_b;
  wire       [7:0]    dSP_525_a;
  wire       [7:0]    dSP_525_d;
  wire       [7:0]    dSP_525_b;
  wire       [7:0]    dSP_526_a;
  wire       [7:0]    dSP_526_d;
  wire       [7:0]    dSP_526_b;
  wire       [7:0]    dSP_527_a;
  wire       [7:0]    dSP_527_d;
  wire       [7:0]    dSP_527_b;
  wire       [7:0]    dSP_528_a;
  wire       [7:0]    dSP_528_d;
  wire       [7:0]    dSP_528_b;
  wire       [7:0]    dSP_529_a;
  wire       [7:0]    dSP_529_d;
  wire       [7:0]    dSP_529_b;
  wire       [7:0]    dSP_530_a;
  wire       [7:0]    dSP_530_d;
  wire       [7:0]    dSP_530_b;
  wire       [7:0]    dSP_531_a;
  wire       [7:0]    dSP_531_d;
  wire       [7:0]    dSP_531_b;
  wire       [7:0]    dSP_532_a;
  wire       [7:0]    dSP_532_d;
  wire       [7:0]    dSP_532_b;
  wire       [7:0]    dSP_533_a;
  wire       [7:0]    dSP_533_d;
  wire       [7:0]    dSP_533_b;
  wire       [7:0]    dSP_534_a;
  wire       [7:0]    dSP_534_d;
  wire       [7:0]    dSP_534_b;
  wire       [7:0]    dSP_535_a;
  wire       [7:0]    dSP_535_d;
  wire       [7:0]    dSP_535_b;
  wire       [7:0]    dSP_536_a;
  wire       [7:0]    dSP_536_d;
  wire       [7:0]    dSP_536_b;
  wire       [7:0]    dSP_537_a;
  wire       [7:0]    dSP_537_d;
  wire       [7:0]    dSP_537_b;
  wire       [7:0]    dSP_538_a;
  wire       [7:0]    dSP_538_d;
  wire       [7:0]    dSP_538_b;
  wire       [7:0]    dSP_539_a;
  wire       [7:0]    dSP_539_d;
  wire       [7:0]    dSP_539_b;
  wire       [7:0]    dSP_540_a;
  wire       [7:0]    dSP_540_d;
  wire       [7:0]    dSP_540_b;
  wire       [7:0]    dSP_541_a;
  wire       [7:0]    dSP_541_d;
  wire       [7:0]    dSP_541_b;
  wire       [7:0]    dSP_542_a;
  wire       [7:0]    dSP_542_d;
  wire       [7:0]    dSP_542_b;
  wire       [7:0]    dSP_543_a;
  wire       [7:0]    dSP_543_d;
  wire       [7:0]    dSP_543_b;
  wire       [7:0]    dSP_544_a;
  wire       [7:0]    dSP_544_d;
  wire       [7:0]    dSP_544_b;
  wire       [7:0]    dSP_545_a;
  wire       [7:0]    dSP_545_d;
  wire       [7:0]    dSP_545_b;
  wire       [7:0]    dSP_546_a;
  wire       [7:0]    dSP_546_d;
  wire       [7:0]    dSP_546_b;
  wire       [7:0]    dSP_547_a;
  wire       [7:0]    dSP_547_d;
  wire       [7:0]    dSP_547_b;
  wire       [7:0]    dSP_548_a;
  wire       [7:0]    dSP_548_d;
  wire       [7:0]    dSP_548_b;
  wire       [7:0]    dSP_549_a;
  wire       [7:0]    dSP_549_d;
  wire       [7:0]    dSP_549_b;
  wire       [7:0]    dSP_550_a;
  wire       [7:0]    dSP_550_d;
  wire       [7:0]    dSP_550_b;
  wire       [7:0]    dSP_551_a;
  wire       [7:0]    dSP_551_d;
  wire       [7:0]    dSP_551_b;
  wire       [7:0]    dSP_552_a;
  wire       [7:0]    dSP_552_d;
  wire       [7:0]    dSP_552_b;
  wire       [7:0]    dSP_553_a;
  wire       [7:0]    dSP_553_d;
  wire       [7:0]    dSP_553_b;
  wire       [7:0]    dSP_554_a;
  wire       [7:0]    dSP_554_d;
  wire       [7:0]    dSP_554_b;
  wire       [7:0]    dSP_555_a;
  wire       [7:0]    dSP_555_d;
  wire       [7:0]    dSP_555_b;
  wire       [7:0]    dSP_556_a;
  wire       [7:0]    dSP_556_d;
  wire       [7:0]    dSP_556_b;
  wire       [7:0]    dSP_557_a;
  wire       [7:0]    dSP_557_d;
  wire       [7:0]    dSP_557_b;
  wire       [7:0]    dSP_558_a;
  wire       [7:0]    dSP_558_d;
  wire       [7:0]    dSP_558_b;
  wire       [7:0]    dSP_559_a;
  wire       [7:0]    dSP_559_d;
  wire       [7:0]    dSP_559_b;
  wire       [7:0]    dSP_560_a;
  wire       [7:0]    dSP_560_d;
  wire       [7:0]    dSP_560_b;
  wire       [7:0]    dSP_561_a;
  wire       [7:0]    dSP_561_d;
  wire       [7:0]    dSP_561_b;
  wire       [7:0]    dSP_562_a;
  wire       [7:0]    dSP_562_d;
  wire       [7:0]    dSP_562_b;
  wire       [7:0]    dSP_563_a;
  wire       [7:0]    dSP_563_d;
  wire       [7:0]    dSP_563_b;
  wire       [7:0]    dSP_564_a;
  wire       [7:0]    dSP_564_d;
  wire       [7:0]    dSP_564_b;
  wire       [7:0]    dSP_565_a;
  wire       [7:0]    dSP_565_d;
  wire       [7:0]    dSP_565_b;
  wire       [7:0]    dSP_566_a;
  wire       [7:0]    dSP_566_d;
  wire       [7:0]    dSP_566_b;
  wire       [7:0]    dSP_567_a;
  wire       [7:0]    dSP_567_d;
  wire       [7:0]    dSP_567_b;
  wire       [7:0]    dSP_568_a;
  wire       [7:0]    dSP_568_d;
  wire       [7:0]    dSP_568_b;
  wire       [7:0]    dSP_569_a;
  wire       [7:0]    dSP_569_d;
  wire       [7:0]    dSP_569_b;
  wire       [7:0]    dSP_570_a;
  wire       [7:0]    dSP_570_d;
  wire       [7:0]    dSP_570_b;
  wire       [7:0]    dSP_571_a;
  wire       [7:0]    dSP_571_d;
  wire       [7:0]    dSP_571_b;
  wire       [7:0]    dSP_572_a;
  wire       [7:0]    dSP_572_d;
  wire       [7:0]    dSP_572_b;
  wire       [7:0]    dSP_573_a;
  wire       [7:0]    dSP_573_d;
  wire       [7:0]    dSP_573_b;
  wire       [7:0]    dSP_574_a;
  wire       [7:0]    dSP_574_d;
  wire       [7:0]    dSP_574_b;
  wire       [7:0]    dSP_575_a;
  wire       [7:0]    dSP_575_d;
  wire       [7:0]    dSP_575_b;
  wire       [7:0]    dSP_576_a;
  wire       [7:0]    dSP_576_d;
  wire       [7:0]    dSP_576_b;
  wire       [7:0]    dSP_577_a;
  wire       [7:0]    dSP_577_d;
  wire       [7:0]    dSP_577_b;
  wire       [7:0]    dSP_578_a;
  wire       [7:0]    dSP_578_d;
  wire       [7:0]    dSP_578_b;
  wire       [7:0]    dSP_579_a;
  wire       [7:0]    dSP_579_d;
  wire       [7:0]    dSP_579_b;
  wire       [7:0]    dSP_580_a;
  wire       [7:0]    dSP_580_d;
  wire       [7:0]    dSP_580_b;
  wire       [7:0]    dSP_581_a;
  wire       [7:0]    dSP_581_d;
  wire       [7:0]    dSP_581_b;
  wire       [7:0]    dSP_582_a;
  wire       [7:0]    dSP_582_d;
  wire       [7:0]    dSP_582_b;
  wire       [7:0]    dSP_583_a;
  wire       [7:0]    dSP_583_d;
  wire       [7:0]    dSP_583_b;
  wire       [7:0]    dSP_584_a;
  wire       [7:0]    dSP_584_d;
  wire       [7:0]    dSP_584_b;
  wire       [7:0]    dSP_585_a;
  wire       [7:0]    dSP_585_d;
  wire       [7:0]    dSP_585_b;
  wire       [7:0]    dSP_586_a;
  wire       [7:0]    dSP_586_d;
  wire       [7:0]    dSP_586_b;
  wire       [7:0]    dSP_587_a;
  wire       [7:0]    dSP_587_d;
  wire       [7:0]    dSP_587_b;
  wire       [7:0]    dSP_588_a;
  wire       [7:0]    dSP_588_d;
  wire       [7:0]    dSP_588_b;
  wire       [7:0]    dSP_589_a;
  wire       [7:0]    dSP_589_d;
  wire       [7:0]    dSP_589_b;
  wire       [7:0]    dSP_590_a;
  wire       [7:0]    dSP_590_d;
  wire       [7:0]    dSP_590_b;
  wire       [7:0]    dSP_591_a;
  wire       [7:0]    dSP_591_d;
  wire       [7:0]    dSP_591_b;
  wire       [7:0]    dSP_592_a;
  wire       [7:0]    dSP_592_d;
  wire       [7:0]    dSP_592_b;
  wire       [7:0]    dSP_593_a;
  wire       [7:0]    dSP_593_d;
  wire       [7:0]    dSP_593_b;
  wire       [7:0]    dSP_594_a;
  wire       [7:0]    dSP_594_d;
  wire       [7:0]    dSP_594_b;
  wire       [7:0]    dSP_595_a;
  wire       [7:0]    dSP_595_d;
  wire       [7:0]    dSP_595_b;
  wire       [7:0]    dSP_596_a;
  wire       [7:0]    dSP_596_d;
  wire       [7:0]    dSP_596_b;
  wire       [7:0]    dSP_597_a;
  wire       [7:0]    dSP_597_d;
  wire       [7:0]    dSP_597_b;
  wire       [7:0]    dSP_598_a;
  wire       [7:0]    dSP_598_d;
  wire       [7:0]    dSP_598_b;
  wire       [7:0]    dSP_599_a;
  wire       [7:0]    dSP_599_d;
  wire       [7:0]    dSP_599_b;
  wire       [7:0]    dSP_600_a;
  wire       [7:0]    dSP_600_d;
  wire       [7:0]    dSP_600_b;
  wire       [7:0]    dSP_601_a;
  wire       [7:0]    dSP_601_d;
  wire       [7:0]    dSP_601_b;
  wire       [7:0]    dSP_602_a;
  wire       [7:0]    dSP_602_d;
  wire       [7:0]    dSP_602_b;
  wire       [7:0]    dSP_603_a;
  wire       [7:0]    dSP_603_d;
  wire       [7:0]    dSP_603_b;
  wire       [7:0]    dSP_604_a;
  wire       [7:0]    dSP_604_d;
  wire       [7:0]    dSP_604_b;
  wire       [7:0]    dSP_605_a;
  wire       [7:0]    dSP_605_d;
  wire       [7:0]    dSP_605_b;
  wire       [7:0]    dSP_606_a;
  wire       [7:0]    dSP_606_d;
  wire       [7:0]    dSP_606_b;
  wire       [7:0]    dSP_607_a;
  wire       [7:0]    dSP_607_d;
  wire       [7:0]    dSP_607_b;
  wire       [7:0]    dSP_608_a;
  wire       [7:0]    dSP_608_d;
  wire       [7:0]    dSP_608_b;
  wire       [7:0]    dSP_609_a;
  wire       [7:0]    dSP_609_d;
  wire       [7:0]    dSP_609_b;
  wire       [7:0]    dSP_610_a;
  wire       [7:0]    dSP_610_d;
  wire       [7:0]    dSP_610_b;
  wire       [7:0]    dSP_611_a;
  wire       [7:0]    dSP_611_d;
  wire       [7:0]    dSP_611_b;
  wire       [7:0]    dSP_612_a;
  wire       [7:0]    dSP_612_d;
  wire       [7:0]    dSP_612_b;
  wire       [7:0]    dSP_613_a;
  wire       [7:0]    dSP_613_d;
  wire       [7:0]    dSP_613_b;
  wire       [7:0]    dSP_614_a;
  wire       [7:0]    dSP_614_d;
  wire       [7:0]    dSP_614_b;
  wire       [7:0]    dSP_615_a;
  wire       [7:0]    dSP_615_d;
  wire       [7:0]    dSP_615_b;
  wire       [7:0]    dSP_616_a;
  wire       [7:0]    dSP_616_d;
  wire       [7:0]    dSP_616_b;
  wire       [7:0]    dSP_617_a;
  wire       [7:0]    dSP_617_d;
  wire       [7:0]    dSP_617_b;
  wire       [7:0]    dSP_618_a;
  wire       [7:0]    dSP_618_d;
  wire       [7:0]    dSP_618_b;
  wire       [7:0]    dSP_619_a;
  wire       [7:0]    dSP_619_d;
  wire       [7:0]    dSP_619_b;
  wire       [7:0]    dSP_620_a;
  wire       [7:0]    dSP_620_d;
  wire       [7:0]    dSP_620_b;
  wire       [7:0]    dSP_621_a;
  wire       [7:0]    dSP_621_d;
  wire       [7:0]    dSP_621_b;
  wire       [7:0]    dSP_622_a;
  wire       [7:0]    dSP_622_d;
  wire       [7:0]    dSP_622_b;
  wire       [7:0]    dSP_623_a;
  wire       [7:0]    dSP_623_d;
  wire       [7:0]    dSP_623_b;
  wire       [7:0]    dSP_624_a;
  wire       [7:0]    dSP_624_d;
  wire       [7:0]    dSP_624_b;
  wire       [7:0]    dSP_625_a;
  wire       [7:0]    dSP_625_d;
  wire       [7:0]    dSP_625_b;
  wire       [7:0]    dSP_626_a;
  wire       [7:0]    dSP_626_d;
  wire       [7:0]    dSP_626_b;
  wire       [7:0]    dSP_627_a;
  wire       [7:0]    dSP_627_d;
  wire       [7:0]    dSP_627_b;
  wire       [7:0]    dSP_628_a;
  wire       [7:0]    dSP_628_d;
  wire       [7:0]    dSP_628_b;
  wire       [7:0]    dSP_629_a;
  wire       [7:0]    dSP_629_d;
  wire       [7:0]    dSP_629_b;
  wire       [7:0]    dSP_630_a;
  wire       [7:0]    dSP_630_d;
  wire       [7:0]    dSP_630_b;
  wire       [7:0]    dSP_631_a;
  wire       [7:0]    dSP_631_d;
  wire       [7:0]    dSP_631_b;
  wire       [7:0]    dSP_632_a;
  wire       [7:0]    dSP_632_d;
  wire       [7:0]    dSP_632_b;
  wire       [7:0]    dSP_633_a;
  wire       [7:0]    dSP_633_d;
  wire       [7:0]    dSP_633_b;
  wire       [7:0]    dSP_634_a;
  wire       [7:0]    dSP_634_d;
  wire       [7:0]    dSP_634_b;
  wire       [7:0]    dSP_635_a;
  wire       [7:0]    dSP_635_d;
  wire       [7:0]    dSP_635_b;
  wire       [7:0]    dSP_636_a;
  wire       [7:0]    dSP_636_d;
  wire       [7:0]    dSP_636_b;
  wire       [7:0]    dSP_637_a;
  wire       [7:0]    dSP_637_d;
  wire       [7:0]    dSP_637_b;
  wire       [7:0]    dSP_638_a;
  wire       [7:0]    dSP_638_d;
  wire       [7:0]    dSP_638_b;
  wire       [7:0]    dSP_639_a;
  wire       [7:0]    dSP_639_d;
  wire       [7:0]    dSP_639_b;
  wire       [7:0]    dSP_640_a;
  wire       [7:0]    dSP_640_d;
  wire       [7:0]    dSP_640_b;
  wire       [7:0]    dSP_641_a;
  wire       [7:0]    dSP_641_d;
  wire       [7:0]    dSP_641_b;
  wire       [7:0]    dSP_642_a;
  wire       [7:0]    dSP_642_d;
  wire       [7:0]    dSP_642_b;
  wire       [7:0]    dSP_643_a;
  wire       [7:0]    dSP_643_d;
  wire       [7:0]    dSP_643_b;
  wire       [7:0]    dSP_644_a;
  wire       [7:0]    dSP_644_d;
  wire       [7:0]    dSP_644_b;
  wire       [7:0]    dSP_645_a;
  wire       [7:0]    dSP_645_d;
  wire       [7:0]    dSP_645_b;
  wire       [7:0]    dSP_646_a;
  wire       [7:0]    dSP_646_d;
  wire       [7:0]    dSP_646_b;
  wire       [7:0]    dSP_647_a;
  wire       [7:0]    dSP_647_d;
  wire       [7:0]    dSP_647_b;
  wire       [7:0]    dSP_648_a;
  wire       [7:0]    dSP_648_d;
  wire       [7:0]    dSP_648_b;
  wire       [7:0]    dSP_649_a;
  wire       [7:0]    dSP_649_d;
  wire       [7:0]    dSP_649_b;
  wire       [7:0]    dSP_650_a;
  wire       [7:0]    dSP_650_d;
  wire       [7:0]    dSP_650_b;
  wire       [7:0]    dSP_651_a;
  wire       [7:0]    dSP_651_d;
  wire       [7:0]    dSP_651_b;
  wire       [7:0]    dSP_652_a;
  wire       [7:0]    dSP_652_d;
  wire       [7:0]    dSP_652_b;
  wire       [7:0]    dSP_653_a;
  wire       [7:0]    dSP_653_d;
  wire       [7:0]    dSP_653_b;
  wire       [7:0]    dSP_654_a;
  wire       [7:0]    dSP_654_d;
  wire       [7:0]    dSP_654_b;
  wire       [7:0]    dSP_655_a;
  wire       [7:0]    dSP_655_d;
  wire       [7:0]    dSP_655_b;
  wire       [7:0]    dSP_656_a;
  wire       [7:0]    dSP_656_d;
  wire       [7:0]    dSP_656_b;
  wire       [7:0]    dSP_657_a;
  wire       [7:0]    dSP_657_d;
  wire       [7:0]    dSP_657_b;
  wire       [7:0]    dSP_658_a;
  wire       [7:0]    dSP_658_d;
  wire       [7:0]    dSP_658_b;
  wire       [7:0]    dSP_659_a;
  wire       [7:0]    dSP_659_d;
  wire       [7:0]    dSP_659_b;
  wire       [7:0]    dSP_660_a;
  wire       [7:0]    dSP_660_d;
  wire       [7:0]    dSP_660_b;
  wire       [7:0]    dSP_661_a;
  wire       [7:0]    dSP_661_d;
  wire       [7:0]    dSP_661_b;
  wire       [7:0]    dSP_662_a;
  wire       [7:0]    dSP_662_d;
  wire       [7:0]    dSP_662_b;
  wire       [7:0]    dSP_663_a;
  wire       [7:0]    dSP_663_d;
  wire       [7:0]    dSP_663_b;
  wire       [7:0]    dSP_664_a;
  wire       [7:0]    dSP_664_d;
  wire       [7:0]    dSP_664_b;
  wire       [7:0]    dSP_665_a;
  wire       [7:0]    dSP_665_d;
  wire       [7:0]    dSP_665_b;
  wire       [7:0]    dSP_666_a;
  wire       [7:0]    dSP_666_d;
  wire       [7:0]    dSP_666_b;
  wire       [7:0]    dSP_667_a;
  wire       [7:0]    dSP_667_d;
  wire       [7:0]    dSP_667_b;
  wire       [7:0]    dSP_668_a;
  wire       [7:0]    dSP_668_d;
  wire       [7:0]    dSP_668_b;
  wire       [7:0]    dSP_669_a;
  wire       [7:0]    dSP_669_d;
  wire       [7:0]    dSP_669_b;
  wire       [7:0]    dSP_670_a;
  wire       [7:0]    dSP_670_d;
  wire       [7:0]    dSP_670_b;
  wire       [7:0]    dSP_671_a;
  wire       [7:0]    dSP_671_d;
  wire       [7:0]    dSP_671_b;
  wire       [7:0]    dSP_672_a;
  wire       [7:0]    dSP_672_d;
  wire       [7:0]    dSP_672_b;
  wire       [7:0]    dSP_673_a;
  wire       [7:0]    dSP_673_d;
  wire       [7:0]    dSP_673_b;
  wire       [7:0]    dSP_674_a;
  wire       [7:0]    dSP_674_d;
  wire       [7:0]    dSP_674_b;
  wire       [7:0]    dSP_675_a;
  wire       [7:0]    dSP_675_d;
  wire       [7:0]    dSP_675_b;
  wire       [7:0]    dSP_676_a;
  wire       [7:0]    dSP_676_d;
  wire       [7:0]    dSP_676_b;
  wire       [7:0]    dSP_677_a;
  wire       [7:0]    dSP_677_d;
  wire       [7:0]    dSP_677_b;
  wire       [7:0]    dSP_678_a;
  wire       [7:0]    dSP_678_d;
  wire       [7:0]    dSP_678_b;
  wire       [7:0]    dSP_679_a;
  wire       [7:0]    dSP_679_d;
  wire       [7:0]    dSP_679_b;
  wire       [7:0]    dSP_680_a;
  wire       [7:0]    dSP_680_d;
  wire       [7:0]    dSP_680_b;
  wire       [7:0]    dSP_681_a;
  wire       [7:0]    dSP_681_d;
  wire       [7:0]    dSP_681_b;
  wire       [7:0]    dSP_682_a;
  wire       [7:0]    dSP_682_d;
  wire       [7:0]    dSP_682_b;
  wire       [7:0]    dSP_683_a;
  wire       [7:0]    dSP_683_d;
  wire       [7:0]    dSP_683_b;
  wire       [7:0]    dSP_684_a;
  wire       [7:0]    dSP_684_d;
  wire       [7:0]    dSP_684_b;
  wire       [7:0]    dSP_685_a;
  wire       [7:0]    dSP_685_d;
  wire       [7:0]    dSP_685_b;
  wire       [7:0]    dSP_686_a;
  wire       [7:0]    dSP_686_d;
  wire       [7:0]    dSP_686_b;
  wire       [7:0]    dSP_687_a;
  wire       [7:0]    dSP_687_d;
  wire       [7:0]    dSP_687_b;
  wire       [7:0]    dSP_688_a;
  wire       [7:0]    dSP_688_d;
  wire       [7:0]    dSP_688_b;
  wire       [7:0]    dSP_689_a;
  wire       [7:0]    dSP_689_d;
  wire       [7:0]    dSP_689_b;
  wire       [7:0]    dSP_690_a;
  wire       [7:0]    dSP_690_d;
  wire       [7:0]    dSP_690_b;
  wire       [7:0]    dSP_691_a;
  wire       [7:0]    dSP_691_d;
  wire       [7:0]    dSP_691_b;
  wire       [7:0]    dSP_692_a;
  wire       [7:0]    dSP_692_d;
  wire       [7:0]    dSP_692_b;
  wire       [7:0]    dSP_693_a;
  wire       [7:0]    dSP_693_d;
  wire       [7:0]    dSP_693_b;
  wire       [7:0]    dSP_694_a;
  wire       [7:0]    dSP_694_d;
  wire       [7:0]    dSP_694_b;
  wire       [7:0]    dSP_695_a;
  wire       [7:0]    dSP_695_d;
  wire       [7:0]    dSP_695_b;
  wire       [7:0]    dSP_696_a;
  wire       [7:0]    dSP_696_d;
  wire       [7:0]    dSP_696_b;
  wire       [7:0]    dSP_697_a;
  wire       [7:0]    dSP_697_d;
  wire       [7:0]    dSP_697_b;
  wire       [7:0]    dSP_698_a;
  wire       [7:0]    dSP_698_d;
  wire       [7:0]    dSP_698_b;
  wire       [7:0]    dSP_699_a;
  wire       [7:0]    dSP_699_d;
  wire       [7:0]    dSP_699_b;
  wire       [7:0]    dSP_700_a;
  wire       [7:0]    dSP_700_d;
  wire       [7:0]    dSP_700_b;
  wire       [7:0]    dSP_701_a;
  wire       [7:0]    dSP_701_d;
  wire       [7:0]    dSP_701_b;
  wire       [7:0]    dSP_702_a;
  wire       [7:0]    dSP_702_d;
  wire       [7:0]    dSP_702_b;
  wire       [7:0]    dSP_703_a;
  wire       [7:0]    dSP_703_d;
  wire       [7:0]    dSP_703_b;
  wire       [7:0]    dSP_704_a;
  wire       [7:0]    dSP_704_d;
  wire       [7:0]    dSP_704_b;
  wire       [7:0]    dSP_705_a;
  wire       [7:0]    dSP_705_d;
  wire       [7:0]    dSP_705_b;
  wire       [7:0]    dSP_706_a;
  wire       [7:0]    dSP_706_d;
  wire       [7:0]    dSP_706_b;
  wire       [7:0]    dSP_707_a;
  wire       [7:0]    dSP_707_d;
  wire       [7:0]    dSP_707_b;
  wire       [7:0]    dSP_708_a;
  wire       [7:0]    dSP_708_d;
  wire       [7:0]    dSP_708_b;
  wire       [7:0]    dSP_709_a;
  wire       [7:0]    dSP_709_d;
  wire       [7:0]    dSP_709_b;
  wire       [7:0]    dSP_710_a;
  wire       [7:0]    dSP_710_d;
  wire       [7:0]    dSP_710_b;
  wire       [7:0]    dSP_711_a;
  wire       [7:0]    dSP_711_d;
  wire       [7:0]    dSP_711_b;
  wire       [7:0]    dSP_712_a;
  wire       [7:0]    dSP_712_d;
  wire       [7:0]    dSP_712_b;
  wire       [7:0]    dSP_713_a;
  wire       [7:0]    dSP_713_d;
  wire       [7:0]    dSP_713_b;
  wire       [7:0]    dSP_714_a;
  wire       [7:0]    dSP_714_d;
  wire       [7:0]    dSP_714_b;
  wire       [7:0]    dSP_715_a;
  wire       [7:0]    dSP_715_d;
  wire       [7:0]    dSP_715_b;
  wire       [7:0]    dSP_716_a;
  wire       [7:0]    dSP_716_d;
  wire       [7:0]    dSP_716_b;
  wire       [7:0]    dSP_717_a;
  wire       [7:0]    dSP_717_d;
  wire       [7:0]    dSP_717_b;
  wire       [7:0]    dSP_718_a;
  wire       [7:0]    dSP_718_d;
  wire       [7:0]    dSP_718_b;
  wire       [7:0]    dSP_719_a;
  wire       [7:0]    dSP_719_d;
  wire       [7:0]    dSP_719_b;
  wire       [7:0]    dSP_720_a;
  wire       [7:0]    dSP_720_d;
  wire       [7:0]    dSP_720_b;
  wire       [7:0]    dSP_721_a;
  wire       [7:0]    dSP_721_d;
  wire       [7:0]    dSP_721_b;
  wire       [7:0]    dSP_722_a;
  wire       [7:0]    dSP_722_d;
  wire       [7:0]    dSP_722_b;
  wire       [7:0]    dSP_723_a;
  wire       [7:0]    dSP_723_d;
  wire       [7:0]    dSP_723_b;
  wire       [7:0]    dSP_724_a;
  wire       [7:0]    dSP_724_d;
  wire       [7:0]    dSP_724_b;
  wire       [7:0]    dSP_725_a;
  wire       [7:0]    dSP_725_d;
  wire       [7:0]    dSP_725_b;
  wire       [7:0]    dSP_726_a;
  wire       [7:0]    dSP_726_d;
  wire       [7:0]    dSP_726_b;
  wire       [7:0]    dSP_727_a;
  wire       [7:0]    dSP_727_d;
  wire       [7:0]    dSP_727_b;
  wire       [7:0]    dSP_728_a;
  wire       [7:0]    dSP_728_d;
  wire       [7:0]    dSP_728_b;
  wire       [7:0]    dSP_729_a;
  wire       [7:0]    dSP_729_d;
  wire       [7:0]    dSP_729_b;
  wire       [7:0]    dSP_730_a;
  wire       [7:0]    dSP_730_d;
  wire       [7:0]    dSP_730_b;
  wire       [7:0]    dSP_731_a;
  wire       [7:0]    dSP_731_d;
  wire       [7:0]    dSP_731_b;
  wire       [7:0]    dSP_732_a;
  wire       [7:0]    dSP_732_d;
  wire       [7:0]    dSP_732_b;
  wire       [7:0]    dSP_733_a;
  wire       [7:0]    dSP_733_d;
  wire       [7:0]    dSP_733_b;
  wire       [7:0]    dSP_734_a;
  wire       [7:0]    dSP_734_d;
  wire       [7:0]    dSP_734_b;
  wire       [7:0]    dSP_735_a;
  wire       [7:0]    dSP_735_d;
  wire       [7:0]    dSP_735_b;
  wire       [7:0]    dSP_736_a;
  wire       [7:0]    dSP_736_d;
  wire       [7:0]    dSP_736_b;
  wire       [7:0]    dSP_737_a;
  wire       [7:0]    dSP_737_d;
  wire       [7:0]    dSP_737_b;
  wire       [7:0]    dSP_738_a;
  wire       [7:0]    dSP_738_d;
  wire       [7:0]    dSP_738_b;
  wire       [7:0]    dSP_739_a;
  wire       [7:0]    dSP_739_d;
  wire       [7:0]    dSP_739_b;
  wire       [7:0]    dSP_740_a;
  wire       [7:0]    dSP_740_d;
  wire       [7:0]    dSP_740_b;
  wire       [7:0]    dSP_741_a;
  wire       [7:0]    dSP_741_d;
  wire       [7:0]    dSP_741_b;
  wire       [7:0]    dSP_742_a;
  wire       [7:0]    dSP_742_d;
  wire       [7:0]    dSP_742_b;
  wire       [7:0]    dSP_743_a;
  wire       [7:0]    dSP_743_d;
  wire       [7:0]    dSP_743_b;
  wire       [7:0]    dSP_744_a;
  wire       [7:0]    dSP_744_d;
  wire       [7:0]    dSP_744_b;
  wire       [7:0]    dSP_745_a;
  wire       [7:0]    dSP_745_d;
  wire       [7:0]    dSP_745_b;
  wire       [7:0]    dSP_746_a;
  wire       [7:0]    dSP_746_d;
  wire       [7:0]    dSP_746_b;
  wire       [7:0]    dSP_747_a;
  wire       [7:0]    dSP_747_d;
  wire       [7:0]    dSP_747_b;
  wire       [7:0]    dSP_748_a;
  wire       [7:0]    dSP_748_d;
  wire       [7:0]    dSP_748_b;
  wire       [7:0]    dSP_749_a;
  wire       [7:0]    dSP_749_d;
  wire       [7:0]    dSP_749_b;
  wire       [7:0]    dSP_750_a;
  wire       [7:0]    dSP_750_d;
  wire       [7:0]    dSP_750_b;
  wire       [7:0]    dSP_751_a;
  wire       [7:0]    dSP_751_d;
  wire       [7:0]    dSP_751_b;
  wire       [7:0]    dSP_752_a;
  wire       [7:0]    dSP_752_d;
  wire       [7:0]    dSP_752_b;
  wire       [7:0]    dSP_753_a;
  wire       [7:0]    dSP_753_d;
  wire       [7:0]    dSP_753_b;
  wire       [7:0]    dSP_754_a;
  wire       [7:0]    dSP_754_d;
  wire       [7:0]    dSP_754_b;
  wire       [7:0]    dSP_755_a;
  wire       [7:0]    dSP_755_d;
  wire       [7:0]    dSP_755_b;
  wire       [7:0]    dSP_756_a;
  wire       [7:0]    dSP_756_d;
  wire       [7:0]    dSP_756_b;
  wire       [7:0]    dSP_757_a;
  wire       [7:0]    dSP_757_d;
  wire       [7:0]    dSP_757_b;
  wire       [7:0]    dSP_758_a;
  wire       [7:0]    dSP_758_d;
  wire       [7:0]    dSP_758_b;
  wire       [7:0]    dSP_759_a;
  wire       [7:0]    dSP_759_d;
  wire       [7:0]    dSP_759_b;
  wire       [7:0]    dSP_760_a;
  wire       [7:0]    dSP_760_d;
  wire       [7:0]    dSP_760_b;
  wire       [7:0]    dSP_761_a;
  wire       [7:0]    dSP_761_d;
  wire       [7:0]    dSP_761_b;
  wire       [7:0]    dSP_762_a;
  wire       [7:0]    dSP_762_d;
  wire       [7:0]    dSP_762_b;
  wire       [7:0]    dSP_763_a;
  wire       [7:0]    dSP_763_d;
  wire       [7:0]    dSP_763_b;
  wire       [7:0]    dSP_764_a;
  wire       [7:0]    dSP_764_d;
  wire       [7:0]    dSP_764_b;
  wire       [7:0]    dSP_765_a;
  wire       [7:0]    dSP_765_d;
  wire       [7:0]    dSP_765_b;
  wire       [7:0]    dSP_766_a;
  wire       [7:0]    dSP_766_d;
  wire       [7:0]    dSP_766_b;
  wire       [7:0]    dSP_767_a;
  wire       [7:0]    dSP_767_d;
  wire       [7:0]    dSP_767_b;
  wire       [7:0]    dSP_768_a;
  wire       [7:0]    dSP_768_d;
  wire       [7:0]    dSP_768_b;
  wire       [7:0]    dSP_769_a;
  wire       [7:0]    dSP_769_d;
  wire       [7:0]    dSP_769_b;
  wire       [7:0]    dSP_770_a;
  wire       [7:0]    dSP_770_d;
  wire       [7:0]    dSP_770_b;
  wire       [7:0]    dSP_771_a;
  wire       [7:0]    dSP_771_d;
  wire       [7:0]    dSP_771_b;
  wire       [7:0]    dSP_772_a;
  wire       [7:0]    dSP_772_d;
  wire       [7:0]    dSP_772_b;
  wire       [7:0]    dSP_773_a;
  wire       [7:0]    dSP_773_d;
  wire       [7:0]    dSP_773_b;
  wire       [7:0]    dSP_774_a;
  wire       [7:0]    dSP_774_d;
  wire       [7:0]    dSP_774_b;
  wire       [7:0]    dSP_775_a;
  wire       [7:0]    dSP_775_d;
  wire       [7:0]    dSP_775_b;
  wire       [7:0]    dSP_776_a;
  wire       [7:0]    dSP_776_d;
  wire       [7:0]    dSP_776_b;
  wire       [7:0]    dSP_777_a;
  wire       [7:0]    dSP_777_d;
  wire       [7:0]    dSP_777_b;
  wire       [7:0]    dSP_778_a;
  wire       [7:0]    dSP_778_d;
  wire       [7:0]    dSP_778_b;
  wire       [7:0]    dSP_779_a;
  wire       [7:0]    dSP_779_d;
  wire       [7:0]    dSP_779_b;
  wire       [7:0]    dSP_780_a;
  wire       [7:0]    dSP_780_d;
  wire       [7:0]    dSP_780_b;
  wire       [7:0]    dSP_781_a;
  wire       [7:0]    dSP_781_d;
  wire       [7:0]    dSP_781_b;
  wire       [7:0]    dSP_782_a;
  wire       [7:0]    dSP_782_d;
  wire       [7:0]    dSP_782_b;
  wire       [7:0]    dSP_783_a;
  wire       [7:0]    dSP_783_d;
  wire       [7:0]    dSP_783_b;
  wire       [7:0]    dSP_784_a;
  wire       [7:0]    dSP_784_d;
  wire       [7:0]    dSP_784_b;
  wire       [7:0]    dSP_785_a;
  wire       [7:0]    dSP_785_d;
  wire       [7:0]    dSP_785_b;
  wire       [7:0]    dSP_786_a;
  wire       [7:0]    dSP_786_d;
  wire       [7:0]    dSP_786_b;
  wire       [7:0]    dSP_787_a;
  wire       [7:0]    dSP_787_d;
  wire       [7:0]    dSP_787_b;
  wire       [7:0]    dSP_788_a;
  wire       [7:0]    dSP_788_d;
  wire       [7:0]    dSP_788_b;
  wire       [7:0]    dSP_789_a;
  wire       [7:0]    dSP_789_d;
  wire       [7:0]    dSP_789_b;
  wire       [7:0]    dSP_790_a;
  wire       [7:0]    dSP_790_d;
  wire       [7:0]    dSP_790_b;
  wire       [7:0]    dSP_791_a;
  wire       [7:0]    dSP_791_d;
  wire       [7:0]    dSP_791_b;
  wire       [7:0]    dSP_792_a;
  wire       [7:0]    dSP_792_d;
  wire       [7:0]    dSP_792_b;
  wire       [7:0]    dSP_793_a;
  wire       [7:0]    dSP_793_d;
  wire       [7:0]    dSP_793_b;
  wire       [7:0]    dSP_794_a;
  wire       [7:0]    dSP_794_d;
  wire       [7:0]    dSP_794_b;
  wire       [7:0]    dSP_795_a;
  wire       [7:0]    dSP_795_d;
  wire       [7:0]    dSP_795_b;
  wire       [7:0]    dSP_796_a;
  wire       [7:0]    dSP_796_d;
  wire       [7:0]    dSP_796_b;
  wire       [7:0]    dSP_797_a;
  wire       [7:0]    dSP_797_d;
  wire       [7:0]    dSP_797_b;
  wire       [7:0]    dSP_798_a;
  wire       [7:0]    dSP_798_d;
  wire       [7:0]    dSP_798_b;
  wire       [7:0]    dSP_799_a;
  wire       [7:0]    dSP_799_d;
  wire       [7:0]    dSP_799_b;
  wire       [7:0]    dSP_800_a;
  wire       [7:0]    dSP_800_d;
  wire       [7:0]    dSP_800_b;
  wire       [7:0]    dSP_801_a;
  wire       [7:0]    dSP_801_d;
  wire       [7:0]    dSP_801_b;
  wire       [7:0]    dSP_802_a;
  wire       [7:0]    dSP_802_d;
  wire       [7:0]    dSP_802_b;
  wire       [7:0]    dSP_803_a;
  wire       [7:0]    dSP_803_d;
  wire       [7:0]    dSP_803_b;
  wire       [7:0]    dSP_804_a;
  wire       [7:0]    dSP_804_d;
  wire       [7:0]    dSP_804_b;
  wire       [7:0]    dSP_805_a;
  wire       [7:0]    dSP_805_d;
  wire       [7:0]    dSP_805_b;
  wire       [7:0]    dSP_806_a;
  wire       [7:0]    dSP_806_d;
  wire       [7:0]    dSP_806_b;
  wire       [7:0]    dSP_807_a;
  wire       [7:0]    dSP_807_d;
  wire       [7:0]    dSP_807_b;
  wire       [7:0]    dSP_808_a;
  wire       [7:0]    dSP_808_d;
  wire       [7:0]    dSP_808_b;
  wire       [7:0]    dSP_809_a;
  wire       [7:0]    dSP_809_d;
  wire       [7:0]    dSP_809_b;
  wire       [7:0]    dSP_810_a;
  wire       [7:0]    dSP_810_d;
  wire       [7:0]    dSP_810_b;
  wire       [7:0]    dSP_811_a;
  wire       [7:0]    dSP_811_d;
  wire       [7:0]    dSP_811_b;
  wire       [7:0]    dSP_812_a;
  wire       [7:0]    dSP_812_d;
  wire       [7:0]    dSP_812_b;
  wire       [7:0]    dSP_813_a;
  wire       [7:0]    dSP_813_d;
  wire       [7:0]    dSP_813_b;
  wire       [7:0]    dSP_814_a;
  wire       [7:0]    dSP_814_d;
  wire       [7:0]    dSP_814_b;
  wire       [7:0]    dSP_815_a;
  wire       [7:0]    dSP_815_d;
  wire       [7:0]    dSP_815_b;
  wire       [7:0]    dSP_816_a;
  wire       [7:0]    dSP_816_d;
  wire       [7:0]    dSP_816_b;
  wire       [7:0]    dSP_817_a;
  wire       [7:0]    dSP_817_d;
  wire       [7:0]    dSP_817_b;
  wire       [7:0]    dSP_818_a;
  wire       [7:0]    dSP_818_d;
  wire       [7:0]    dSP_818_b;
  wire       [7:0]    dSP_819_a;
  wire       [7:0]    dSP_819_d;
  wire       [7:0]    dSP_819_b;
  wire       [7:0]    dSP_820_a;
  wire       [7:0]    dSP_820_d;
  wire       [7:0]    dSP_820_b;
  wire       [7:0]    dSP_821_a;
  wire       [7:0]    dSP_821_d;
  wire       [7:0]    dSP_821_b;
  wire       [7:0]    dSP_822_a;
  wire       [7:0]    dSP_822_d;
  wire       [7:0]    dSP_822_b;
  wire       [7:0]    dSP_823_a;
  wire       [7:0]    dSP_823_d;
  wire       [7:0]    dSP_823_b;
  wire       [7:0]    dSP_824_a;
  wire       [7:0]    dSP_824_d;
  wire       [7:0]    dSP_824_b;
  wire       [7:0]    dSP_825_a;
  wire       [7:0]    dSP_825_d;
  wire       [7:0]    dSP_825_b;
  wire       [7:0]    dSP_826_a;
  wire       [7:0]    dSP_826_d;
  wire       [7:0]    dSP_826_b;
  wire       [7:0]    dSP_827_a;
  wire       [7:0]    dSP_827_d;
  wire       [7:0]    dSP_827_b;
  wire       [7:0]    dSP_828_a;
  wire       [7:0]    dSP_828_d;
  wire       [7:0]    dSP_828_b;
  wire       [7:0]    dSP_829_a;
  wire       [7:0]    dSP_829_d;
  wire       [7:0]    dSP_829_b;
  wire       [7:0]    dSP_830_a;
  wire       [7:0]    dSP_830_d;
  wire       [7:0]    dSP_830_b;
  wire       [7:0]    dSP_831_a;
  wire       [7:0]    dSP_831_d;
  wire       [7:0]    dSP_831_b;
  wire       [7:0]    dSP_832_a;
  wire       [7:0]    dSP_832_d;
  wire       [7:0]    dSP_832_b;
  wire       [7:0]    dSP_833_a;
  wire       [7:0]    dSP_833_d;
  wire       [7:0]    dSP_833_b;
  wire       [7:0]    dSP_834_a;
  wire       [7:0]    dSP_834_d;
  wire       [7:0]    dSP_834_b;
  wire       [7:0]    dSP_835_a;
  wire       [7:0]    dSP_835_d;
  wire       [7:0]    dSP_835_b;
  wire       [7:0]    dSP_836_a;
  wire       [7:0]    dSP_836_d;
  wire       [7:0]    dSP_836_b;
  wire       [7:0]    dSP_837_a;
  wire       [7:0]    dSP_837_d;
  wire       [7:0]    dSP_837_b;
  wire       [7:0]    dSP_838_a;
  wire       [7:0]    dSP_838_d;
  wire       [7:0]    dSP_838_b;
  wire       [7:0]    dSP_839_a;
  wire       [7:0]    dSP_839_d;
  wire       [7:0]    dSP_839_b;
  wire       [7:0]    dSP_840_a;
  wire       [7:0]    dSP_840_d;
  wire       [7:0]    dSP_840_b;
  wire       [7:0]    dSP_841_a;
  wire       [7:0]    dSP_841_d;
  wire       [7:0]    dSP_841_b;
  wire       [7:0]    dSP_842_a;
  wire       [7:0]    dSP_842_d;
  wire       [7:0]    dSP_842_b;
  wire       [7:0]    dSP_843_a;
  wire       [7:0]    dSP_843_d;
  wire       [7:0]    dSP_843_b;
  wire       [7:0]    dSP_844_a;
  wire       [7:0]    dSP_844_d;
  wire       [7:0]    dSP_844_b;
  wire       [7:0]    dSP_845_a;
  wire       [7:0]    dSP_845_d;
  wire       [7:0]    dSP_845_b;
  wire       [7:0]    dSP_846_a;
  wire       [7:0]    dSP_846_d;
  wire       [7:0]    dSP_846_b;
  wire       [7:0]    dSP_847_a;
  wire       [7:0]    dSP_847_d;
  wire       [7:0]    dSP_847_b;
  wire       [7:0]    dSP_848_a;
  wire       [7:0]    dSP_848_d;
  wire       [7:0]    dSP_848_b;
  wire       [7:0]    dSP_849_a;
  wire       [7:0]    dSP_849_d;
  wire       [7:0]    dSP_849_b;
  wire       [7:0]    dSP_850_a;
  wire       [7:0]    dSP_850_d;
  wire       [7:0]    dSP_850_b;
  wire       [7:0]    dSP_851_a;
  wire       [7:0]    dSP_851_d;
  wire       [7:0]    dSP_851_b;
  wire       [7:0]    dSP_852_a;
  wire       [7:0]    dSP_852_d;
  wire       [7:0]    dSP_852_b;
  wire       [7:0]    dSP_853_a;
  wire       [7:0]    dSP_853_d;
  wire       [7:0]    dSP_853_b;
  wire       [7:0]    dSP_854_a;
  wire       [7:0]    dSP_854_d;
  wire       [7:0]    dSP_854_b;
  wire       [7:0]    dSP_855_a;
  wire       [7:0]    dSP_855_d;
  wire       [7:0]    dSP_855_b;
  wire       [7:0]    dSP_856_a;
  wire       [7:0]    dSP_856_d;
  wire       [7:0]    dSP_856_b;
  wire       [7:0]    dSP_857_a;
  wire       [7:0]    dSP_857_d;
  wire       [7:0]    dSP_857_b;
  wire       [7:0]    dSP_858_a;
  wire       [7:0]    dSP_858_d;
  wire       [7:0]    dSP_858_b;
  wire       [7:0]    dSP_859_a;
  wire       [7:0]    dSP_859_d;
  wire       [7:0]    dSP_859_b;
  wire       [7:0]    dSP_860_a;
  wire       [7:0]    dSP_860_d;
  wire       [7:0]    dSP_860_b;
  wire       [7:0]    dSP_861_a;
  wire       [7:0]    dSP_861_d;
  wire       [7:0]    dSP_861_b;
  wire       [7:0]    dSP_862_a;
  wire       [7:0]    dSP_862_d;
  wire       [7:0]    dSP_862_b;
  wire       [7:0]    dSP_863_a;
  wire       [7:0]    dSP_863_d;
  wire       [7:0]    dSP_863_b;
  wire       [7:0]    dSP_864_a;
  wire       [7:0]    dSP_864_d;
  wire       [7:0]    dSP_864_b;
  wire       [7:0]    dSP_865_a;
  wire       [7:0]    dSP_865_d;
  wire       [7:0]    dSP_865_b;
  wire       [7:0]    dSP_866_a;
  wire       [7:0]    dSP_866_d;
  wire       [7:0]    dSP_866_b;
  wire       [7:0]    dSP_867_a;
  wire       [7:0]    dSP_867_d;
  wire       [7:0]    dSP_867_b;
  wire       [7:0]    dSP_868_a;
  wire       [7:0]    dSP_868_d;
  wire       [7:0]    dSP_868_b;
  wire       [7:0]    dSP_869_a;
  wire       [7:0]    dSP_869_d;
  wire       [7:0]    dSP_869_b;
  wire       [7:0]    dSP_870_a;
  wire       [7:0]    dSP_870_d;
  wire       [7:0]    dSP_870_b;
  wire       [7:0]    dSP_871_a;
  wire       [7:0]    dSP_871_d;
  wire       [7:0]    dSP_871_b;
  wire       [7:0]    dSP_872_a;
  wire       [7:0]    dSP_872_d;
  wire       [7:0]    dSP_872_b;
  wire       [7:0]    dSP_873_a;
  wire       [7:0]    dSP_873_d;
  wire       [7:0]    dSP_873_b;
  wire       [7:0]    dSP_874_a;
  wire       [7:0]    dSP_874_d;
  wire       [7:0]    dSP_874_b;
  wire       [7:0]    dSP_875_a;
  wire       [7:0]    dSP_875_d;
  wire       [7:0]    dSP_875_b;
  wire       [7:0]    dSP_876_a;
  wire       [7:0]    dSP_876_d;
  wire       [7:0]    dSP_876_b;
  wire       [7:0]    dSP_877_a;
  wire       [7:0]    dSP_877_d;
  wire       [7:0]    dSP_877_b;
  wire       [7:0]    dSP_878_a;
  wire       [7:0]    dSP_878_d;
  wire       [7:0]    dSP_878_b;
  wire       [7:0]    dSP_879_a;
  wire       [7:0]    dSP_879_d;
  wire       [7:0]    dSP_879_b;
  wire       [7:0]    dSP_880_a;
  wire       [7:0]    dSP_880_d;
  wire       [7:0]    dSP_880_b;
  wire       [7:0]    dSP_881_a;
  wire       [7:0]    dSP_881_d;
  wire       [7:0]    dSP_881_b;
  wire       [7:0]    dSP_882_a;
  wire       [7:0]    dSP_882_d;
  wire       [7:0]    dSP_882_b;
  wire       [7:0]    dSP_883_a;
  wire       [7:0]    dSP_883_d;
  wire       [7:0]    dSP_883_b;
  wire       [7:0]    dSP_884_a;
  wire       [7:0]    dSP_884_d;
  wire       [7:0]    dSP_884_b;
  wire       [7:0]    dSP_885_a;
  wire       [7:0]    dSP_885_d;
  wire       [7:0]    dSP_885_b;
  wire       [7:0]    dSP_886_a;
  wire       [7:0]    dSP_886_d;
  wire       [7:0]    dSP_886_b;
  wire       [7:0]    dSP_887_a;
  wire       [7:0]    dSP_887_d;
  wire       [7:0]    dSP_887_b;
  wire       [7:0]    dSP_888_a;
  wire       [7:0]    dSP_888_d;
  wire       [7:0]    dSP_888_b;
  wire       [7:0]    dSP_889_a;
  wire       [7:0]    dSP_889_d;
  wire       [7:0]    dSP_889_b;
  wire       [7:0]    dSP_890_a;
  wire       [7:0]    dSP_890_d;
  wire       [7:0]    dSP_890_b;
  wire       [7:0]    dSP_891_a;
  wire       [7:0]    dSP_891_d;
  wire       [7:0]    dSP_891_b;
  wire       [7:0]    dSP_892_a;
  wire       [7:0]    dSP_892_d;
  wire       [7:0]    dSP_892_b;
  wire       [7:0]    dSP_893_a;
  wire       [7:0]    dSP_893_d;
  wire       [7:0]    dSP_893_b;
  wire       [7:0]    dSP_894_a;
  wire       [7:0]    dSP_894_d;
  wire       [7:0]    dSP_894_b;
  wire       [7:0]    dSP_895_a;
  wire       [7:0]    dSP_895_d;
  wire       [7:0]    dSP_895_b;
  wire       [7:0]    dSP_896_a;
  wire       [7:0]    dSP_896_d;
  wire       [7:0]    dSP_896_b;
  wire       [7:0]    dSP_897_a;
  wire       [7:0]    dSP_897_d;
  wire       [7:0]    dSP_897_b;
  wire       [7:0]    dSP_898_a;
  wire       [7:0]    dSP_898_d;
  wire       [7:0]    dSP_898_b;
  wire       [7:0]    dSP_899_a;
  wire       [7:0]    dSP_899_d;
  wire       [7:0]    dSP_899_b;
  wire       [7:0]    dSP_900_a;
  wire       [7:0]    dSP_900_d;
  wire       [7:0]    dSP_900_b;
  wire       [7:0]    dSP_901_a;
  wire       [7:0]    dSP_901_d;
  wire       [7:0]    dSP_901_b;
  wire       [7:0]    dSP_902_a;
  wire       [7:0]    dSP_902_d;
  wire       [7:0]    dSP_902_b;
  wire       [7:0]    dSP_903_a;
  wire       [7:0]    dSP_903_d;
  wire       [7:0]    dSP_903_b;
  wire       [7:0]    dSP_904_a;
  wire       [7:0]    dSP_904_d;
  wire       [7:0]    dSP_904_b;
  wire       [7:0]    dSP_905_a;
  wire       [7:0]    dSP_905_d;
  wire       [7:0]    dSP_905_b;
  wire       [7:0]    dSP_906_a;
  wire       [7:0]    dSP_906_d;
  wire       [7:0]    dSP_906_b;
  wire       [7:0]    dSP_907_a;
  wire       [7:0]    dSP_907_d;
  wire       [7:0]    dSP_907_b;
  wire       [7:0]    dSP_908_a;
  wire       [7:0]    dSP_908_d;
  wire       [7:0]    dSP_908_b;
  wire       [7:0]    dSP_909_a;
  wire       [7:0]    dSP_909_d;
  wire       [7:0]    dSP_909_b;
  wire       [7:0]    dSP_910_a;
  wire       [7:0]    dSP_910_d;
  wire       [7:0]    dSP_910_b;
  wire       [7:0]    dSP_911_a;
  wire       [7:0]    dSP_911_d;
  wire       [7:0]    dSP_911_b;
  wire       [7:0]    dSP_912_a;
  wire       [7:0]    dSP_912_d;
  wire       [7:0]    dSP_912_b;
  wire       [7:0]    dSP_913_a;
  wire       [7:0]    dSP_913_d;
  wire       [7:0]    dSP_913_b;
  wire       [7:0]    dSP_914_a;
  wire       [7:0]    dSP_914_d;
  wire       [7:0]    dSP_914_b;
  wire       [7:0]    dSP_915_a;
  wire       [7:0]    dSP_915_d;
  wire       [7:0]    dSP_915_b;
  wire       [7:0]    dSP_916_a;
  wire       [7:0]    dSP_916_d;
  wire       [7:0]    dSP_916_b;
  wire       [7:0]    dSP_917_a;
  wire       [7:0]    dSP_917_d;
  wire       [7:0]    dSP_917_b;
  wire       [7:0]    dSP_918_a;
  wire       [7:0]    dSP_918_d;
  wire       [7:0]    dSP_918_b;
  wire       [7:0]    dSP_919_a;
  wire       [7:0]    dSP_919_d;
  wire       [7:0]    dSP_919_b;
  wire       [7:0]    dSP_920_a;
  wire       [7:0]    dSP_920_d;
  wire       [7:0]    dSP_920_b;
  wire       [7:0]    dSP_921_a;
  wire       [7:0]    dSP_921_d;
  wire       [7:0]    dSP_921_b;
  wire       [7:0]    dSP_922_a;
  wire       [7:0]    dSP_922_d;
  wire       [7:0]    dSP_922_b;
  wire       [7:0]    dSP_923_a;
  wire       [7:0]    dSP_923_d;
  wire       [7:0]    dSP_923_b;
  wire       [7:0]    dSP_924_a;
  wire       [7:0]    dSP_924_d;
  wire       [7:0]    dSP_924_b;
  wire       [7:0]    dSP_925_a;
  wire       [7:0]    dSP_925_d;
  wire       [7:0]    dSP_925_b;
  wire       [7:0]    dSP_926_a;
  wire       [7:0]    dSP_926_d;
  wire       [7:0]    dSP_926_b;
  wire       [7:0]    dSP_927_a;
  wire       [7:0]    dSP_927_d;
  wire       [7:0]    dSP_927_b;
  wire       [7:0]    dSP_928_a;
  wire       [7:0]    dSP_928_d;
  wire       [7:0]    dSP_928_b;
  wire       [7:0]    dSP_929_a;
  wire       [7:0]    dSP_929_d;
  wire       [7:0]    dSP_929_b;
  wire       [7:0]    dSP_930_a;
  wire       [7:0]    dSP_930_d;
  wire       [7:0]    dSP_930_b;
  wire       [7:0]    dSP_931_a;
  wire       [7:0]    dSP_931_d;
  wire       [7:0]    dSP_931_b;
  wire       [7:0]    dSP_932_a;
  wire       [7:0]    dSP_932_d;
  wire       [7:0]    dSP_932_b;
  wire       [7:0]    dSP_933_a;
  wire       [7:0]    dSP_933_d;
  wire       [7:0]    dSP_933_b;
  wire       [7:0]    dSP_934_a;
  wire       [7:0]    dSP_934_d;
  wire       [7:0]    dSP_934_b;
  wire       [7:0]    dSP_935_a;
  wire       [7:0]    dSP_935_d;
  wire       [7:0]    dSP_935_b;
  wire       [7:0]    dSP_936_a;
  wire       [7:0]    dSP_936_d;
  wire       [7:0]    dSP_936_b;
  wire       [7:0]    dSP_937_a;
  wire       [7:0]    dSP_937_d;
  wire       [7:0]    dSP_937_b;
  wire       [7:0]    dSP_938_a;
  wire       [7:0]    dSP_938_d;
  wire       [7:0]    dSP_938_b;
  wire       [7:0]    dSP_939_a;
  wire       [7:0]    dSP_939_d;
  wire       [7:0]    dSP_939_b;
  wire       [7:0]    dSP_940_a;
  wire       [7:0]    dSP_940_d;
  wire       [7:0]    dSP_940_b;
  wire       [7:0]    dSP_941_a;
  wire       [7:0]    dSP_941_d;
  wire       [7:0]    dSP_941_b;
  wire       [7:0]    dSP_942_a;
  wire       [7:0]    dSP_942_d;
  wire       [7:0]    dSP_942_b;
  wire       [7:0]    dSP_943_a;
  wire       [7:0]    dSP_943_d;
  wire       [7:0]    dSP_943_b;
  wire       [7:0]    dSP_944_a;
  wire       [7:0]    dSP_944_d;
  wire       [7:0]    dSP_944_b;
  wire       [7:0]    dSP_945_a;
  wire       [7:0]    dSP_945_d;
  wire       [7:0]    dSP_945_b;
  wire       [7:0]    dSP_946_a;
  wire       [7:0]    dSP_946_d;
  wire       [7:0]    dSP_946_b;
  wire       [7:0]    dSP_947_a;
  wire       [7:0]    dSP_947_d;
  wire       [7:0]    dSP_947_b;
  wire       [7:0]    dSP_948_a;
  wire       [7:0]    dSP_948_d;
  wire       [7:0]    dSP_948_b;
  wire       [7:0]    dSP_949_a;
  wire       [7:0]    dSP_949_d;
  wire       [7:0]    dSP_949_b;
  wire       [7:0]    dSP_950_a;
  wire       [7:0]    dSP_950_d;
  wire       [7:0]    dSP_950_b;
  wire       [7:0]    dSP_951_a;
  wire       [7:0]    dSP_951_d;
  wire       [7:0]    dSP_951_b;
  wire       [7:0]    dSP_952_a;
  wire       [7:0]    dSP_952_d;
  wire       [7:0]    dSP_952_b;
  wire       [7:0]    dSP_953_a;
  wire       [7:0]    dSP_953_d;
  wire       [7:0]    dSP_953_b;
  wire       [7:0]    dSP_954_a;
  wire       [7:0]    dSP_954_d;
  wire       [7:0]    dSP_954_b;
  wire       [7:0]    dSP_955_a;
  wire       [7:0]    dSP_955_d;
  wire       [7:0]    dSP_955_b;
  wire       [7:0]    dSP_956_a;
  wire       [7:0]    dSP_956_d;
  wire       [7:0]    dSP_956_b;
  wire       [7:0]    dSP_957_a;
  wire       [7:0]    dSP_957_d;
  wire       [7:0]    dSP_957_b;
  wire       [7:0]    dSP_958_a;
  wire       [7:0]    dSP_958_d;
  wire       [7:0]    dSP_958_b;
  wire       [7:0]    dSP_959_a;
  wire       [7:0]    dSP_959_d;
  wire       [7:0]    dSP_959_b;
  wire       [7:0]    dSP_960_a;
  wire       [7:0]    dSP_960_d;
  wire       [7:0]    dSP_960_b;
  wire       [7:0]    dSP_961_a;
  wire       [7:0]    dSP_961_d;
  wire       [7:0]    dSP_961_b;
  wire       [7:0]    dSP_962_a;
  wire       [7:0]    dSP_962_d;
  wire       [7:0]    dSP_962_b;
  wire       [7:0]    dSP_963_a;
  wire       [7:0]    dSP_963_d;
  wire       [7:0]    dSP_963_b;
  wire       [7:0]    dSP_964_a;
  wire       [7:0]    dSP_964_d;
  wire       [7:0]    dSP_964_b;
  wire       [7:0]    dSP_965_a;
  wire       [7:0]    dSP_965_d;
  wire       [7:0]    dSP_965_b;
  wire       [7:0]    dSP_966_a;
  wire       [7:0]    dSP_966_d;
  wire       [7:0]    dSP_966_b;
  wire       [7:0]    dSP_967_a;
  wire       [7:0]    dSP_967_d;
  wire       [7:0]    dSP_967_b;
  wire       [7:0]    dSP_968_a;
  wire       [7:0]    dSP_968_d;
  wire       [7:0]    dSP_968_b;
  wire       [7:0]    dSP_969_a;
  wire       [7:0]    dSP_969_d;
  wire       [7:0]    dSP_969_b;
  wire       [7:0]    dSP_970_a;
  wire       [7:0]    dSP_970_d;
  wire       [7:0]    dSP_970_b;
  wire       [7:0]    dSP_971_a;
  wire       [7:0]    dSP_971_d;
  wire       [7:0]    dSP_971_b;
  wire       [7:0]    dSP_972_a;
  wire       [7:0]    dSP_972_d;
  wire       [7:0]    dSP_972_b;
  wire       [7:0]    dSP_973_a;
  wire       [7:0]    dSP_973_d;
  wire       [7:0]    dSP_973_b;
  wire       [7:0]    dSP_974_a;
  wire       [7:0]    dSP_974_d;
  wire       [7:0]    dSP_974_b;
  wire       [7:0]    dSP_975_a;
  wire       [7:0]    dSP_975_d;
  wire       [7:0]    dSP_975_b;
  wire       [7:0]    dSP_976_a;
  wire       [7:0]    dSP_976_d;
  wire       [7:0]    dSP_976_b;
  wire       [7:0]    dSP_977_a;
  wire       [7:0]    dSP_977_d;
  wire       [7:0]    dSP_977_b;
  wire       [7:0]    dSP_978_a;
  wire       [7:0]    dSP_978_d;
  wire       [7:0]    dSP_978_b;
  wire       [7:0]    dSP_979_a;
  wire       [7:0]    dSP_979_d;
  wire       [7:0]    dSP_979_b;
  wire       [7:0]    dSP_980_a;
  wire       [7:0]    dSP_980_d;
  wire       [7:0]    dSP_980_b;
  wire       [7:0]    dSP_981_a;
  wire       [7:0]    dSP_981_d;
  wire       [7:0]    dSP_981_b;
  wire       [7:0]    dSP_982_a;
  wire       [7:0]    dSP_982_d;
  wire       [7:0]    dSP_982_b;
  wire       [7:0]    dSP_983_a;
  wire       [7:0]    dSP_983_d;
  wire       [7:0]    dSP_983_b;
  wire       [7:0]    dSP_984_a;
  wire       [7:0]    dSP_984_d;
  wire       [7:0]    dSP_984_b;
  wire       [7:0]    dSP_985_a;
  wire       [7:0]    dSP_985_d;
  wire       [7:0]    dSP_985_b;
  wire       [7:0]    dSP_986_a;
  wire       [7:0]    dSP_986_d;
  wire       [7:0]    dSP_986_b;
  wire       [7:0]    dSP_987_a;
  wire       [7:0]    dSP_987_d;
  wire       [7:0]    dSP_987_b;
  wire       [7:0]    dSP_988_a;
  wire       [7:0]    dSP_988_d;
  wire       [7:0]    dSP_988_b;
  wire       [7:0]    dSP_989_a;
  wire       [7:0]    dSP_989_d;
  wire       [7:0]    dSP_989_b;
  wire       [7:0]    dSP_990_a;
  wire       [7:0]    dSP_990_d;
  wire       [7:0]    dSP_990_b;
  wire       [7:0]    dSP_991_a;
  wire       [7:0]    dSP_991_d;
  wire       [7:0]    dSP_991_b;
  wire       [7:0]    dSP_992_a;
  wire       [7:0]    dSP_992_d;
  wire       [7:0]    dSP_992_b;
  wire       [7:0]    dSP_993_a;
  wire       [7:0]    dSP_993_d;
  wire       [7:0]    dSP_993_b;
  wire       [7:0]    dSP_994_a;
  wire       [7:0]    dSP_994_d;
  wire       [7:0]    dSP_994_b;
  wire       [7:0]    dSP_995_a;
  wire       [7:0]    dSP_995_d;
  wire       [7:0]    dSP_995_b;
  wire       [7:0]    dSP_996_a;
  wire       [7:0]    dSP_996_d;
  wire       [7:0]    dSP_996_b;
  wire       [7:0]    dSP_997_a;
  wire       [7:0]    dSP_997_d;
  wire       [7:0]    dSP_997_b;
  wire       [7:0]    dSP_998_a;
  wire       [7:0]    dSP_998_d;
  wire       [7:0]    dSP_998_b;
  wire       [7:0]    dSP_999_a;
  wire       [7:0]    dSP_999_d;
  wire       [7:0]    dSP_999_b;
  wire       [7:0]    dSP_1000_a;
  wire       [7:0]    dSP_1000_d;
  wire       [7:0]    dSP_1000_b;
  wire       [7:0]    dSP_1001_a;
  wire       [7:0]    dSP_1001_d;
  wire       [7:0]    dSP_1001_b;
  wire       [7:0]    dSP_1002_a;
  wire       [7:0]    dSP_1002_d;
  wire       [7:0]    dSP_1002_b;
  wire       [7:0]    dSP_1003_a;
  wire       [7:0]    dSP_1003_d;
  wire       [7:0]    dSP_1003_b;
  wire       [7:0]    dSP_1004_a;
  wire       [7:0]    dSP_1004_d;
  wire       [7:0]    dSP_1004_b;
  wire       [7:0]    dSP_1005_a;
  wire       [7:0]    dSP_1005_d;
  wire       [7:0]    dSP_1005_b;
  wire       [7:0]    dSP_1006_a;
  wire       [7:0]    dSP_1006_d;
  wire       [7:0]    dSP_1006_b;
  wire       [7:0]    dSP_1007_a;
  wire       [7:0]    dSP_1007_d;
  wire       [7:0]    dSP_1007_b;
  wire       [7:0]    dSP_1008_a;
  wire       [7:0]    dSP_1008_d;
  wire       [7:0]    dSP_1008_b;
  wire       [7:0]    dSP_1009_a;
  wire       [7:0]    dSP_1009_d;
  wire       [7:0]    dSP_1009_b;
  wire       [7:0]    dSP_1010_a;
  wire       [7:0]    dSP_1010_d;
  wire       [7:0]    dSP_1010_b;
  wire       [7:0]    dSP_1011_a;
  wire       [7:0]    dSP_1011_d;
  wire       [7:0]    dSP_1011_b;
  wire       [7:0]    dSP_1012_a;
  wire       [7:0]    dSP_1012_d;
  wire       [7:0]    dSP_1012_b;
  wire       [7:0]    dSP_1013_a;
  wire       [7:0]    dSP_1013_d;
  wire       [7:0]    dSP_1013_b;
  wire       [7:0]    dSP_1014_a;
  wire       [7:0]    dSP_1014_d;
  wire       [7:0]    dSP_1014_b;
  wire       [7:0]    dSP_1015_a;
  wire       [7:0]    dSP_1015_d;
  wire       [7:0]    dSP_1015_b;
  wire       [7:0]    dSP_1016_a;
  wire       [7:0]    dSP_1016_d;
  wire       [7:0]    dSP_1016_b;
  wire       [7:0]    dSP_1017_a;
  wire       [7:0]    dSP_1017_d;
  wire       [7:0]    dSP_1017_b;
  wire       [7:0]    dSP_1018_a;
  wire       [7:0]    dSP_1018_d;
  wire       [7:0]    dSP_1018_b;
  wire       [7:0]    dSP_1019_a;
  wire       [7:0]    dSP_1019_d;
  wire       [7:0]    dSP_1019_b;
  wire       [7:0]    dSP_1020_a;
  wire       [7:0]    dSP_1020_d;
  wire       [7:0]    dSP_1020_b;
  wire       [7:0]    dSP_1021_a;
  wire       [7:0]    dSP_1021_d;
  wire       [7:0]    dSP_1021_b;
  wire       [7:0]    dSP_1022_a;
  wire       [7:0]    dSP_1022_d;
  wire       [7:0]    dSP_1022_b;
  wire       [7:0]    dSP_1023_a;
  wire       [7:0]    dSP_1023_d;
  wire       [7:0]    dSP_1023_b;
  wire       [7:0]    dSP_1024_a;
  wire       [7:0]    dSP_1024_d;
  wire       [7:0]    dSP_1024_b;
  wire       [7:0]    dSP_1025_a;
  wire       [7:0]    dSP_1025_d;
  wire       [7:0]    dSP_1025_b;
  wire       [7:0]    dSP_1026_a;
  wire       [7:0]    dSP_1026_d;
  wire       [7:0]    dSP_1026_b;
  wire       [7:0]    dSP_1027_a;
  wire       [7:0]    dSP_1027_d;
  wire       [7:0]    dSP_1027_b;
  wire       [7:0]    dSP_1028_a;
  wire       [7:0]    dSP_1028_d;
  wire       [7:0]    dSP_1028_b;
  wire       [7:0]    dSP_1029_a;
  wire       [7:0]    dSP_1029_d;
  wire       [7:0]    dSP_1029_b;
  wire       [7:0]    dSP_1030_a;
  wire       [7:0]    dSP_1030_d;
  wire       [7:0]    dSP_1030_b;
  wire       [7:0]    dSP_1031_a;
  wire       [7:0]    dSP_1031_d;
  wire       [7:0]    dSP_1031_b;
  wire       [7:0]    dSP_1032_a;
  wire       [7:0]    dSP_1032_d;
  wire       [7:0]    dSP_1032_b;
  wire       [7:0]    dSP_1033_a;
  wire       [7:0]    dSP_1033_d;
  wire       [7:0]    dSP_1033_b;
  wire       [7:0]    dSP_1034_a;
  wire       [7:0]    dSP_1034_d;
  wire       [7:0]    dSP_1034_b;
  wire       [7:0]    dSP_1035_a;
  wire       [7:0]    dSP_1035_d;
  wire       [7:0]    dSP_1035_b;
  wire       [7:0]    dSP_1036_a;
  wire       [7:0]    dSP_1036_d;
  wire       [7:0]    dSP_1036_b;
  wire       [7:0]    dSP_1037_a;
  wire       [7:0]    dSP_1037_d;
  wire       [7:0]    dSP_1037_b;
  wire       [7:0]    dSP_1038_a;
  wire       [7:0]    dSP_1038_d;
  wire       [7:0]    dSP_1038_b;
  wire       [7:0]    dSP_1039_a;
  wire       [7:0]    dSP_1039_d;
  wire       [7:0]    dSP_1039_b;
  wire       [7:0]    dSP_1040_a;
  wire       [7:0]    dSP_1040_d;
  wire       [7:0]    dSP_1040_b;
  wire       [7:0]    dSP_1041_a;
  wire       [7:0]    dSP_1041_d;
  wire       [7:0]    dSP_1041_b;
  wire       [7:0]    dSP_1042_a;
  wire       [7:0]    dSP_1042_d;
  wire       [7:0]    dSP_1042_b;
  wire       [7:0]    dSP_1043_a;
  wire       [7:0]    dSP_1043_d;
  wire       [7:0]    dSP_1043_b;
  wire       [7:0]    dSP_1044_a;
  wire       [7:0]    dSP_1044_d;
  wire       [7:0]    dSP_1044_b;
  wire       [7:0]    dSP_1045_a;
  wire       [7:0]    dSP_1045_d;
  wire       [7:0]    dSP_1045_b;
  wire       [7:0]    dSP_1046_a;
  wire       [7:0]    dSP_1046_d;
  wire       [7:0]    dSP_1046_b;
  wire       [7:0]    dSP_1047_a;
  wire       [7:0]    dSP_1047_d;
  wire       [7:0]    dSP_1047_b;
  wire       [7:0]    dSP_1048_a;
  wire       [7:0]    dSP_1048_d;
  wire       [7:0]    dSP_1048_b;
  wire       [7:0]    dSP_1049_a;
  wire       [7:0]    dSP_1049_d;
  wire       [7:0]    dSP_1049_b;
  wire       [7:0]    dSP_1050_a;
  wire       [7:0]    dSP_1050_d;
  wire       [7:0]    dSP_1050_b;
  wire       [7:0]    dSP_1051_a;
  wire       [7:0]    dSP_1051_d;
  wire       [7:0]    dSP_1051_b;
  wire       [7:0]    dSP_1052_a;
  wire       [7:0]    dSP_1052_d;
  wire       [7:0]    dSP_1052_b;
  wire       [7:0]    dSP_1053_a;
  wire       [7:0]    dSP_1053_d;
  wire       [7:0]    dSP_1053_b;
  wire       [7:0]    dSP_1054_a;
  wire       [7:0]    dSP_1054_d;
  wire       [7:0]    dSP_1054_b;
  wire       [7:0]    dSP_1055_a;
  wire       [7:0]    dSP_1055_d;
  wire       [7:0]    dSP_1055_b;
  wire       [7:0]    dSP_1056_a;
  wire       [7:0]    dSP_1056_d;
  wire       [7:0]    dSP_1056_b;
  wire       [7:0]    dSP_1057_a;
  wire       [7:0]    dSP_1057_d;
  wire       [7:0]    dSP_1057_b;
  wire       [7:0]    dSP_1058_a;
  wire       [7:0]    dSP_1058_d;
  wire       [7:0]    dSP_1058_b;
  wire       [7:0]    dSP_1059_a;
  wire       [7:0]    dSP_1059_d;
  wire       [7:0]    dSP_1059_b;
  wire       [7:0]    dSP_1060_a;
  wire       [7:0]    dSP_1060_d;
  wire       [7:0]    dSP_1060_b;
  wire       [7:0]    dSP_1061_a;
  wire       [7:0]    dSP_1061_d;
  wire       [7:0]    dSP_1061_b;
  wire       [7:0]    dSP_1062_a;
  wire       [7:0]    dSP_1062_d;
  wire       [7:0]    dSP_1062_b;
  wire       [7:0]    dSP_1063_a;
  wire       [7:0]    dSP_1063_d;
  wire       [7:0]    dSP_1063_b;
  wire       [7:0]    dSP_1064_a;
  wire       [7:0]    dSP_1064_d;
  wire       [7:0]    dSP_1064_b;
  wire       [7:0]    dSP_1065_a;
  wire       [7:0]    dSP_1065_d;
  wire       [7:0]    dSP_1065_b;
  wire       [7:0]    dSP_1066_a;
  wire       [7:0]    dSP_1066_d;
  wire       [7:0]    dSP_1066_b;
  wire       [7:0]    dSP_1067_a;
  wire       [7:0]    dSP_1067_d;
  wire       [7:0]    dSP_1067_b;
  wire       [7:0]    dSP_1068_a;
  wire       [7:0]    dSP_1068_d;
  wire       [7:0]    dSP_1068_b;
  wire       [7:0]    dSP_1069_a;
  wire       [7:0]    dSP_1069_d;
  wire       [7:0]    dSP_1069_b;
  wire       [7:0]    dSP_1070_a;
  wire       [7:0]    dSP_1070_d;
  wire       [7:0]    dSP_1070_b;
  wire       [7:0]    dSP_1071_a;
  wire       [7:0]    dSP_1071_d;
  wire       [7:0]    dSP_1071_b;
  wire       [7:0]    dSP_1072_a;
  wire       [7:0]    dSP_1072_d;
  wire       [7:0]    dSP_1072_b;
  wire       [7:0]    dSP_1073_a;
  wire       [7:0]    dSP_1073_d;
  wire       [7:0]    dSP_1073_b;
  wire       [7:0]    dSP_1074_a;
  wire       [7:0]    dSP_1074_d;
  wire       [7:0]    dSP_1074_b;
  wire       [7:0]    dSP_1075_a;
  wire       [7:0]    dSP_1075_d;
  wire       [7:0]    dSP_1075_b;
  wire       [7:0]    dSP_1076_a;
  wire       [7:0]    dSP_1076_d;
  wire       [7:0]    dSP_1076_b;
  wire       [7:0]    dSP_1077_a;
  wire       [7:0]    dSP_1077_d;
  wire       [7:0]    dSP_1077_b;
  wire       [7:0]    dSP_1078_a;
  wire       [7:0]    dSP_1078_d;
  wire       [7:0]    dSP_1078_b;
  wire       [7:0]    dSP_1079_a;
  wire       [7:0]    dSP_1079_d;
  wire       [7:0]    dSP_1079_b;
  wire       [7:0]    dSP_1080_a;
  wire       [7:0]    dSP_1080_d;
  wire       [7:0]    dSP_1080_b;
  wire       [7:0]    dSP_1081_a;
  wire       [7:0]    dSP_1081_d;
  wire       [7:0]    dSP_1081_b;
  wire       [7:0]    dSP_1082_a;
  wire       [7:0]    dSP_1082_d;
  wire       [7:0]    dSP_1082_b;
  wire       [7:0]    dSP_1083_a;
  wire       [7:0]    dSP_1083_d;
  wire       [7:0]    dSP_1083_b;
  wire       [7:0]    dSP_1084_a;
  wire       [7:0]    dSP_1084_d;
  wire       [7:0]    dSP_1084_b;
  wire       [7:0]    dSP_1085_a;
  wire       [7:0]    dSP_1085_d;
  wire       [7:0]    dSP_1085_b;
  wire       [7:0]    dSP_1086_a;
  wire       [7:0]    dSP_1086_d;
  wire       [7:0]    dSP_1086_b;
  wire       [7:0]    dSP_1087_a;
  wire       [7:0]    dSP_1087_d;
  wire       [7:0]    dSP_1087_b;
  wire       [7:0]    dSP_1088_a;
  wire       [7:0]    dSP_1088_d;
  wire       [7:0]    dSP_1088_b;
  wire       [7:0]    dSP_1089_a;
  wire       [7:0]    dSP_1089_d;
  wire       [7:0]    dSP_1089_b;
  wire       [7:0]    dSP_1090_a;
  wire       [7:0]    dSP_1090_d;
  wire       [7:0]    dSP_1090_b;
  wire       [7:0]    dSP_1091_a;
  wire       [7:0]    dSP_1091_d;
  wire       [7:0]    dSP_1091_b;
  wire       [7:0]    dSP_1092_a;
  wire       [7:0]    dSP_1092_d;
  wire       [7:0]    dSP_1092_b;
  wire       [7:0]    dSP_1093_a;
  wire       [7:0]    dSP_1093_d;
  wire       [7:0]    dSP_1093_b;
  wire       [7:0]    dSP_1094_a;
  wire       [7:0]    dSP_1094_d;
  wire       [7:0]    dSP_1094_b;
  wire       [7:0]    dSP_1095_a;
  wire       [7:0]    dSP_1095_d;
  wire       [7:0]    dSP_1095_b;
  wire       [7:0]    dSP_1096_a;
  wire       [7:0]    dSP_1096_d;
  wire       [7:0]    dSP_1096_b;
  wire       [7:0]    dSP_1097_a;
  wire       [7:0]    dSP_1097_d;
  wire       [7:0]    dSP_1097_b;
  wire       [7:0]    dSP_1098_a;
  wire       [7:0]    dSP_1098_d;
  wire       [7:0]    dSP_1098_b;
  wire       [7:0]    dSP_1099_a;
  wire       [7:0]    dSP_1099_d;
  wire       [7:0]    dSP_1099_b;
  wire       [7:0]    dSP_1100_a;
  wire       [7:0]    dSP_1100_d;
  wire       [7:0]    dSP_1100_b;
  wire       [7:0]    dSP_1101_a;
  wire       [7:0]    dSP_1101_d;
  wire       [7:0]    dSP_1101_b;
  wire       [7:0]    dSP_1102_a;
  wire       [7:0]    dSP_1102_d;
  wire       [7:0]    dSP_1102_b;
  wire       [7:0]    dSP_1103_a;
  wire       [7:0]    dSP_1103_d;
  wire       [7:0]    dSP_1103_b;
  wire       [7:0]    dSP_1104_a;
  wire       [7:0]    dSP_1104_d;
  wire       [7:0]    dSP_1104_b;
  wire       [7:0]    dSP_1105_a;
  wire       [7:0]    dSP_1105_d;
  wire       [7:0]    dSP_1105_b;
  wire       [7:0]    dSP_1106_a;
  wire       [7:0]    dSP_1106_d;
  wire       [7:0]    dSP_1106_b;
  wire       [7:0]    dSP_1107_a;
  wire       [7:0]    dSP_1107_d;
  wire       [7:0]    dSP_1107_b;
  wire       [7:0]    dSP_1108_a;
  wire       [7:0]    dSP_1108_d;
  wire       [7:0]    dSP_1108_b;
  wire       [7:0]    dSP_1109_a;
  wire       [7:0]    dSP_1109_d;
  wire       [7:0]    dSP_1109_b;
  wire       [7:0]    dSP_1110_a;
  wire       [7:0]    dSP_1110_d;
  wire       [7:0]    dSP_1110_b;
  wire       [7:0]    dSP_1111_a;
  wire       [7:0]    dSP_1111_d;
  wire       [7:0]    dSP_1111_b;
  wire       [7:0]    dSP_1112_a;
  wire       [7:0]    dSP_1112_d;
  wire       [7:0]    dSP_1112_b;
  wire       [7:0]    dSP_1113_a;
  wire       [7:0]    dSP_1113_d;
  wire       [7:0]    dSP_1113_b;
  wire       [7:0]    dSP_1114_a;
  wire       [7:0]    dSP_1114_d;
  wire       [7:0]    dSP_1114_b;
  wire       [7:0]    dSP_1115_a;
  wire       [7:0]    dSP_1115_d;
  wire       [7:0]    dSP_1115_b;
  wire       [7:0]    dSP_1116_a;
  wire       [7:0]    dSP_1116_d;
  wire       [7:0]    dSP_1116_b;
  wire       [7:0]    dSP_1117_a;
  wire       [7:0]    dSP_1117_d;
  wire       [7:0]    dSP_1117_b;
  wire       [7:0]    dSP_1118_a;
  wire       [7:0]    dSP_1118_d;
  wire       [7:0]    dSP_1118_b;
  wire       [7:0]    dSP_1119_a;
  wire       [7:0]    dSP_1119_d;
  wire       [7:0]    dSP_1119_b;
  wire       [7:0]    dSP_1120_a;
  wire       [7:0]    dSP_1120_d;
  wire       [7:0]    dSP_1120_b;
  wire       [7:0]    dSP_1121_a;
  wire       [7:0]    dSP_1121_d;
  wire       [7:0]    dSP_1121_b;
  wire       [7:0]    dSP_1122_a;
  wire       [7:0]    dSP_1122_d;
  wire       [7:0]    dSP_1122_b;
  wire       [7:0]    dSP_1123_a;
  wire       [7:0]    dSP_1123_d;
  wire       [7:0]    dSP_1123_b;
  wire       [7:0]    dSP_1124_a;
  wire       [7:0]    dSP_1124_d;
  wire       [7:0]    dSP_1124_b;
  wire       [7:0]    dSP_1125_a;
  wire       [7:0]    dSP_1125_d;
  wire       [7:0]    dSP_1125_b;
  wire       [7:0]    dSP_1126_a;
  wire       [7:0]    dSP_1126_d;
  wire       [7:0]    dSP_1126_b;
  wire       [7:0]    dSP_1127_a;
  wire       [7:0]    dSP_1127_d;
  wire       [7:0]    dSP_1127_b;
  wire       [7:0]    dSP_1128_a;
  wire       [7:0]    dSP_1128_d;
  wire       [7:0]    dSP_1128_b;
  wire       [7:0]    dSP_1129_a;
  wire       [7:0]    dSP_1129_d;
  wire       [7:0]    dSP_1129_b;
  wire       [7:0]    dSP_1130_a;
  wire       [7:0]    dSP_1130_d;
  wire       [7:0]    dSP_1130_b;
  wire       [7:0]    dSP_1131_a;
  wire       [7:0]    dSP_1131_d;
  wire       [7:0]    dSP_1131_b;
  wire       [7:0]    dSP_1132_a;
  wire       [7:0]    dSP_1132_d;
  wire       [7:0]    dSP_1132_b;
  wire       [7:0]    dSP_1133_a;
  wire       [7:0]    dSP_1133_d;
  wire       [7:0]    dSP_1133_b;
  wire       [7:0]    dSP_1134_a;
  wire       [7:0]    dSP_1134_d;
  wire       [7:0]    dSP_1134_b;
  wire       [7:0]    dSP_1135_a;
  wire       [7:0]    dSP_1135_d;
  wire       [7:0]    dSP_1135_b;
  wire       [7:0]    dSP_1136_a;
  wire       [7:0]    dSP_1136_d;
  wire       [7:0]    dSP_1136_b;
  wire       [7:0]    dSP_1137_a;
  wire       [7:0]    dSP_1137_d;
  wire       [7:0]    dSP_1137_b;
  wire       [7:0]    dSP_1138_a;
  wire       [7:0]    dSP_1138_d;
  wire       [7:0]    dSP_1138_b;
  wire       [7:0]    dSP_1139_a;
  wire       [7:0]    dSP_1139_d;
  wire       [7:0]    dSP_1139_b;
  wire       [7:0]    dSP_1140_a;
  wire       [7:0]    dSP_1140_d;
  wire       [7:0]    dSP_1140_b;
  wire       [7:0]    dSP_1141_a;
  wire       [7:0]    dSP_1141_d;
  wire       [7:0]    dSP_1141_b;
  wire       [7:0]    dSP_1142_a;
  wire       [7:0]    dSP_1142_d;
  wire       [7:0]    dSP_1142_b;
  wire       [7:0]    dSP_1143_a;
  wire       [7:0]    dSP_1143_d;
  wire       [7:0]    dSP_1143_b;
  wire       [7:0]    dSP_1144_a;
  wire       [7:0]    dSP_1144_d;
  wire       [7:0]    dSP_1144_b;
  wire       [7:0]    dSP_1145_a;
  wire       [7:0]    dSP_1145_d;
  wire       [7:0]    dSP_1145_b;
  wire       [7:0]    dSP_1146_a;
  wire       [7:0]    dSP_1146_d;
  wire       [7:0]    dSP_1146_b;
  wire       [7:0]    dSP_1147_a;
  wire       [7:0]    dSP_1147_d;
  wire       [7:0]    dSP_1147_b;
  wire       [7:0]    dSP_1148_a;
  wire       [7:0]    dSP_1148_d;
  wire       [7:0]    dSP_1148_b;
  wire       [7:0]    dSP_1149_a;
  wire       [7:0]    dSP_1149_d;
  wire       [7:0]    dSP_1149_b;
  wire       [7:0]    dSP_1150_a;
  wire       [7:0]    dSP_1150_d;
  wire       [7:0]    dSP_1150_b;
  wire       [7:0]    dSP_1151_a;
  wire       [7:0]    dSP_1151_d;
  wire       [7:0]    dSP_1151_b;
  wire       [7:0]    dSP_1152_a;
  wire       [7:0]    dSP_1152_d;
  wire       [7:0]    dSP_1152_b;
  wire       [31:0]   addKernel_A_0;
  wire       [31:0]   addKernel_A_1;
  wire       [31:0]   addKernel_A_2;
  wire       [31:0]   addKernel_A_3;
  wire       [31:0]   addKernel_A_4;
  wire       [31:0]   addKernel_A_5;
  wire       [31:0]   addKernel_A_6;
  wire       [31:0]   addKernel_A_7;
  wire       [31:0]   addKernel_A_8;
  wire       [31:0]   addKernel_1_A_0;
  wire       [31:0]   addKernel_1_A_1;
  wire       [31:0]   addKernel_1_A_2;
  wire       [31:0]   addKernel_1_A_3;
  wire       [31:0]   addKernel_1_A_4;
  wire       [31:0]   addKernel_1_A_5;
  wire       [31:0]   addKernel_1_A_6;
  wire       [31:0]   addKernel_1_A_7;
  wire       [31:0]   addKernel_1_A_8;
  wire       [31:0]   addKernel_2_A_0;
  wire       [31:0]   addKernel_2_A_1;
  wire       [31:0]   addKernel_2_A_2;
  wire       [31:0]   addKernel_2_A_3;
  wire       [31:0]   addKernel_2_A_4;
  wire       [31:0]   addKernel_2_A_5;
  wire       [31:0]   addKernel_2_A_6;
  wire       [31:0]   addKernel_2_A_7;
  wire       [31:0]   addKernel_2_A_8;
  wire       [31:0]   addKernel_3_A_0;
  wire       [31:0]   addKernel_3_A_1;
  wire       [31:0]   addKernel_3_A_2;
  wire       [31:0]   addKernel_3_A_3;
  wire       [31:0]   addKernel_3_A_4;
  wire       [31:0]   addKernel_3_A_5;
  wire       [31:0]   addKernel_3_A_6;
  wire       [31:0]   addKernel_3_A_7;
  wire       [31:0]   addKernel_3_A_8;
  wire       [31:0]   addKernel_4_A_0;
  wire       [31:0]   addKernel_4_A_1;
  wire       [31:0]   addKernel_4_A_2;
  wire       [31:0]   addKernel_4_A_3;
  wire       [31:0]   addKernel_4_A_4;
  wire       [31:0]   addKernel_4_A_5;
  wire       [31:0]   addKernel_4_A_6;
  wire       [31:0]   addKernel_4_A_7;
  wire       [31:0]   addKernel_4_A_8;
  wire       [31:0]   addKernel_5_A_0;
  wire       [31:0]   addKernel_5_A_1;
  wire       [31:0]   addKernel_5_A_2;
  wire       [31:0]   addKernel_5_A_3;
  wire       [31:0]   addKernel_5_A_4;
  wire       [31:0]   addKernel_5_A_5;
  wire       [31:0]   addKernel_5_A_6;
  wire       [31:0]   addKernel_5_A_7;
  wire       [31:0]   addKernel_5_A_8;
  wire       [31:0]   addKernel_6_A_0;
  wire       [31:0]   addKernel_6_A_1;
  wire       [31:0]   addKernel_6_A_2;
  wire       [31:0]   addKernel_6_A_3;
  wire       [31:0]   addKernel_6_A_4;
  wire       [31:0]   addKernel_6_A_5;
  wire       [31:0]   addKernel_6_A_6;
  wire       [31:0]   addKernel_6_A_7;
  wire       [31:0]   addKernel_6_A_8;
  wire       [31:0]   addKernel_7_A_0;
  wire       [31:0]   addKernel_7_A_1;
  wire       [31:0]   addKernel_7_A_2;
  wire       [31:0]   addKernel_7_A_3;
  wire       [31:0]   addKernel_7_A_4;
  wire       [31:0]   addKernel_7_A_5;
  wire       [31:0]   addKernel_7_A_6;
  wire       [31:0]   addKernel_7_A_7;
  wire       [31:0]   addKernel_7_A_8;
  wire       [31:0]   addKernel_8_A_0;
  wire       [31:0]   addKernel_8_A_1;
  wire       [31:0]   addKernel_8_A_2;
  wire       [31:0]   addKernel_8_A_3;
  wire       [31:0]   addKernel_8_A_4;
  wire       [31:0]   addKernel_8_A_5;
  wire       [31:0]   addKernel_8_A_6;
  wire       [31:0]   addKernel_8_A_7;
  wire       [31:0]   addKernel_8_A_8;
  wire       [31:0]   addKernel_9_A_0;
  wire       [31:0]   addKernel_9_A_1;
  wire       [31:0]   addKernel_9_A_2;
  wire       [31:0]   addKernel_9_A_3;
  wire       [31:0]   addKernel_9_A_4;
  wire       [31:0]   addKernel_9_A_5;
  wire       [31:0]   addKernel_9_A_6;
  wire       [31:0]   addKernel_9_A_7;
  wire       [31:0]   addKernel_9_A_8;
  wire       [31:0]   addKernel_10_A_0;
  wire       [31:0]   addKernel_10_A_1;
  wire       [31:0]   addKernel_10_A_2;
  wire       [31:0]   addKernel_10_A_3;
  wire       [31:0]   addKernel_10_A_4;
  wire       [31:0]   addKernel_10_A_5;
  wire       [31:0]   addKernel_10_A_6;
  wire       [31:0]   addKernel_10_A_7;
  wire       [31:0]   addKernel_10_A_8;
  wire       [31:0]   addKernel_11_A_0;
  wire       [31:0]   addKernel_11_A_1;
  wire       [31:0]   addKernel_11_A_2;
  wire       [31:0]   addKernel_11_A_3;
  wire       [31:0]   addKernel_11_A_4;
  wire       [31:0]   addKernel_11_A_5;
  wire       [31:0]   addKernel_11_A_6;
  wire       [31:0]   addKernel_11_A_7;
  wire       [31:0]   addKernel_11_A_8;
  wire       [31:0]   addKernel_12_A_0;
  wire       [31:0]   addKernel_12_A_1;
  wire       [31:0]   addKernel_12_A_2;
  wire       [31:0]   addKernel_12_A_3;
  wire       [31:0]   addKernel_12_A_4;
  wire       [31:0]   addKernel_12_A_5;
  wire       [31:0]   addKernel_12_A_6;
  wire       [31:0]   addKernel_12_A_7;
  wire       [31:0]   addKernel_12_A_8;
  wire       [31:0]   addKernel_13_A_0;
  wire       [31:0]   addKernel_13_A_1;
  wire       [31:0]   addKernel_13_A_2;
  wire       [31:0]   addKernel_13_A_3;
  wire       [31:0]   addKernel_13_A_4;
  wire       [31:0]   addKernel_13_A_5;
  wire       [31:0]   addKernel_13_A_6;
  wire       [31:0]   addKernel_13_A_7;
  wire       [31:0]   addKernel_13_A_8;
  wire       [31:0]   addKernel_14_A_0;
  wire       [31:0]   addKernel_14_A_1;
  wire       [31:0]   addKernel_14_A_2;
  wire       [31:0]   addKernel_14_A_3;
  wire       [31:0]   addKernel_14_A_4;
  wire       [31:0]   addKernel_14_A_5;
  wire       [31:0]   addKernel_14_A_6;
  wire       [31:0]   addKernel_14_A_7;
  wire       [31:0]   addKernel_14_A_8;
  wire       [31:0]   addKernel_15_A_0;
  wire       [31:0]   addKernel_15_A_1;
  wire       [31:0]   addKernel_15_A_2;
  wire       [31:0]   addKernel_15_A_3;
  wire       [31:0]   addKernel_15_A_4;
  wire       [31:0]   addKernel_15_A_5;
  wire       [31:0]   addKernel_15_A_6;
  wire       [31:0]   addKernel_15_A_7;
  wire       [31:0]   addKernel_15_A_8;
  wire       [31:0]   addKernel_16_A_0;
  wire       [31:0]   addKernel_16_A_1;
  wire       [31:0]   addKernel_16_A_2;
  wire       [31:0]   addKernel_16_A_3;
  wire       [31:0]   addKernel_16_A_4;
  wire       [31:0]   addKernel_16_A_5;
  wire       [31:0]   addKernel_16_A_6;
  wire       [31:0]   addKernel_16_A_7;
  wire       [31:0]   addKernel_16_A_8;
  wire       [31:0]   addKernel_17_A_0;
  wire       [31:0]   addKernel_17_A_1;
  wire       [31:0]   addKernel_17_A_2;
  wire       [31:0]   addKernel_17_A_3;
  wire       [31:0]   addKernel_17_A_4;
  wire       [31:0]   addKernel_17_A_5;
  wire       [31:0]   addKernel_17_A_6;
  wire       [31:0]   addKernel_17_A_7;
  wire       [31:0]   addKernel_17_A_8;
  wire       [31:0]   addKernel_18_A_0;
  wire       [31:0]   addKernel_18_A_1;
  wire       [31:0]   addKernel_18_A_2;
  wire       [31:0]   addKernel_18_A_3;
  wire       [31:0]   addKernel_18_A_4;
  wire       [31:0]   addKernel_18_A_5;
  wire       [31:0]   addKernel_18_A_6;
  wire       [31:0]   addKernel_18_A_7;
  wire       [31:0]   addKernel_18_A_8;
  wire       [31:0]   addKernel_19_A_0;
  wire       [31:0]   addKernel_19_A_1;
  wire       [31:0]   addKernel_19_A_2;
  wire       [31:0]   addKernel_19_A_3;
  wire       [31:0]   addKernel_19_A_4;
  wire       [31:0]   addKernel_19_A_5;
  wire       [31:0]   addKernel_19_A_6;
  wire       [31:0]   addKernel_19_A_7;
  wire       [31:0]   addKernel_19_A_8;
  wire       [31:0]   addKernel_20_A_0;
  wire       [31:0]   addKernel_20_A_1;
  wire       [31:0]   addKernel_20_A_2;
  wire       [31:0]   addKernel_20_A_3;
  wire       [31:0]   addKernel_20_A_4;
  wire       [31:0]   addKernel_20_A_5;
  wire       [31:0]   addKernel_20_A_6;
  wire       [31:0]   addKernel_20_A_7;
  wire       [31:0]   addKernel_20_A_8;
  wire       [31:0]   addKernel_21_A_0;
  wire       [31:0]   addKernel_21_A_1;
  wire       [31:0]   addKernel_21_A_2;
  wire       [31:0]   addKernel_21_A_3;
  wire       [31:0]   addKernel_21_A_4;
  wire       [31:0]   addKernel_21_A_5;
  wire       [31:0]   addKernel_21_A_6;
  wire       [31:0]   addKernel_21_A_7;
  wire       [31:0]   addKernel_21_A_8;
  wire       [31:0]   addKernel_22_A_0;
  wire       [31:0]   addKernel_22_A_1;
  wire       [31:0]   addKernel_22_A_2;
  wire       [31:0]   addKernel_22_A_3;
  wire       [31:0]   addKernel_22_A_4;
  wire       [31:0]   addKernel_22_A_5;
  wire       [31:0]   addKernel_22_A_6;
  wire       [31:0]   addKernel_22_A_7;
  wire       [31:0]   addKernel_22_A_8;
  wire       [31:0]   addKernel_23_A_0;
  wire       [31:0]   addKernel_23_A_1;
  wire       [31:0]   addKernel_23_A_2;
  wire       [31:0]   addKernel_23_A_3;
  wire       [31:0]   addKernel_23_A_4;
  wire       [31:0]   addKernel_23_A_5;
  wire       [31:0]   addKernel_23_A_6;
  wire       [31:0]   addKernel_23_A_7;
  wire       [31:0]   addKernel_23_A_8;
  wire       [31:0]   addKernel_24_A_0;
  wire       [31:0]   addKernel_24_A_1;
  wire       [31:0]   addKernel_24_A_2;
  wire       [31:0]   addKernel_24_A_3;
  wire       [31:0]   addKernel_24_A_4;
  wire       [31:0]   addKernel_24_A_5;
  wire       [31:0]   addKernel_24_A_6;
  wire       [31:0]   addKernel_24_A_7;
  wire       [31:0]   addKernel_24_A_8;
  wire       [31:0]   addKernel_25_A_0;
  wire       [31:0]   addKernel_25_A_1;
  wire       [31:0]   addKernel_25_A_2;
  wire       [31:0]   addKernel_25_A_3;
  wire       [31:0]   addKernel_25_A_4;
  wire       [31:0]   addKernel_25_A_5;
  wire       [31:0]   addKernel_25_A_6;
  wire       [31:0]   addKernel_25_A_7;
  wire       [31:0]   addKernel_25_A_8;
  wire       [31:0]   addKernel_26_A_0;
  wire       [31:0]   addKernel_26_A_1;
  wire       [31:0]   addKernel_26_A_2;
  wire       [31:0]   addKernel_26_A_3;
  wire       [31:0]   addKernel_26_A_4;
  wire       [31:0]   addKernel_26_A_5;
  wire       [31:0]   addKernel_26_A_6;
  wire       [31:0]   addKernel_26_A_7;
  wire       [31:0]   addKernel_26_A_8;
  wire       [31:0]   addKernel_27_A_0;
  wire       [31:0]   addKernel_27_A_1;
  wire       [31:0]   addKernel_27_A_2;
  wire       [31:0]   addKernel_27_A_3;
  wire       [31:0]   addKernel_27_A_4;
  wire       [31:0]   addKernel_27_A_5;
  wire       [31:0]   addKernel_27_A_6;
  wire       [31:0]   addKernel_27_A_7;
  wire       [31:0]   addKernel_27_A_8;
  wire       [31:0]   addKernel_28_A_0;
  wire       [31:0]   addKernel_28_A_1;
  wire       [31:0]   addKernel_28_A_2;
  wire       [31:0]   addKernel_28_A_3;
  wire       [31:0]   addKernel_28_A_4;
  wire       [31:0]   addKernel_28_A_5;
  wire       [31:0]   addKernel_28_A_6;
  wire       [31:0]   addKernel_28_A_7;
  wire       [31:0]   addKernel_28_A_8;
  wire       [31:0]   addKernel_29_A_0;
  wire       [31:0]   addKernel_29_A_1;
  wire       [31:0]   addKernel_29_A_2;
  wire       [31:0]   addKernel_29_A_3;
  wire       [31:0]   addKernel_29_A_4;
  wire       [31:0]   addKernel_29_A_5;
  wire       [31:0]   addKernel_29_A_6;
  wire       [31:0]   addKernel_29_A_7;
  wire       [31:0]   addKernel_29_A_8;
  wire       [31:0]   addKernel_30_A_0;
  wire       [31:0]   addKernel_30_A_1;
  wire       [31:0]   addKernel_30_A_2;
  wire       [31:0]   addKernel_30_A_3;
  wire       [31:0]   addKernel_30_A_4;
  wire       [31:0]   addKernel_30_A_5;
  wire       [31:0]   addKernel_30_A_6;
  wire       [31:0]   addKernel_30_A_7;
  wire       [31:0]   addKernel_30_A_8;
  wire       [31:0]   addKernel_31_A_0;
  wire       [31:0]   addKernel_31_A_1;
  wire       [31:0]   addKernel_31_A_2;
  wire       [31:0]   addKernel_31_A_3;
  wire       [31:0]   addKernel_31_A_4;
  wire       [31:0]   addKernel_31_A_5;
  wire       [31:0]   addKernel_31_A_6;
  wire       [31:0]   addKernel_31_A_7;
  wire       [31:0]   addKernel_31_A_8;
  wire       [31:0]   addKernel_32_A_0;
  wire       [31:0]   addKernel_32_A_1;
  wire       [31:0]   addKernel_32_A_2;
  wire       [31:0]   addKernel_32_A_3;
  wire       [31:0]   addKernel_32_A_4;
  wire       [31:0]   addKernel_32_A_5;
  wire       [31:0]   addKernel_32_A_6;
  wire       [31:0]   addKernel_32_A_7;
  wire       [31:0]   addKernel_32_A_8;
  wire       [31:0]   addKernel_33_A_0;
  wire       [31:0]   addKernel_33_A_1;
  wire       [31:0]   addKernel_33_A_2;
  wire       [31:0]   addKernel_33_A_3;
  wire       [31:0]   addKernel_33_A_4;
  wire       [31:0]   addKernel_33_A_5;
  wire       [31:0]   addKernel_33_A_6;
  wire       [31:0]   addKernel_33_A_7;
  wire       [31:0]   addKernel_33_A_8;
  wire       [31:0]   addKernel_34_A_0;
  wire       [31:0]   addKernel_34_A_1;
  wire       [31:0]   addKernel_34_A_2;
  wire       [31:0]   addKernel_34_A_3;
  wire       [31:0]   addKernel_34_A_4;
  wire       [31:0]   addKernel_34_A_5;
  wire       [31:0]   addKernel_34_A_6;
  wire       [31:0]   addKernel_34_A_7;
  wire       [31:0]   addKernel_34_A_8;
  wire       [31:0]   addKernel_35_A_0;
  wire       [31:0]   addKernel_35_A_1;
  wire       [31:0]   addKernel_35_A_2;
  wire       [31:0]   addKernel_35_A_3;
  wire       [31:0]   addKernel_35_A_4;
  wire       [31:0]   addKernel_35_A_5;
  wire       [31:0]   addKernel_35_A_6;
  wire       [31:0]   addKernel_35_A_7;
  wire       [31:0]   addKernel_35_A_8;
  wire       [31:0]   addKernel_36_A_0;
  wire       [31:0]   addKernel_36_A_1;
  wire       [31:0]   addKernel_36_A_2;
  wire       [31:0]   addKernel_36_A_3;
  wire       [31:0]   addKernel_36_A_4;
  wire       [31:0]   addKernel_36_A_5;
  wire       [31:0]   addKernel_36_A_6;
  wire       [31:0]   addKernel_36_A_7;
  wire       [31:0]   addKernel_36_A_8;
  wire       [31:0]   addKernel_37_A_0;
  wire       [31:0]   addKernel_37_A_1;
  wire       [31:0]   addKernel_37_A_2;
  wire       [31:0]   addKernel_37_A_3;
  wire       [31:0]   addKernel_37_A_4;
  wire       [31:0]   addKernel_37_A_5;
  wire       [31:0]   addKernel_37_A_6;
  wire       [31:0]   addKernel_37_A_7;
  wire       [31:0]   addKernel_37_A_8;
  wire       [31:0]   addKernel_38_A_0;
  wire       [31:0]   addKernel_38_A_1;
  wire       [31:0]   addKernel_38_A_2;
  wire       [31:0]   addKernel_38_A_3;
  wire       [31:0]   addKernel_38_A_4;
  wire       [31:0]   addKernel_38_A_5;
  wire       [31:0]   addKernel_38_A_6;
  wire       [31:0]   addKernel_38_A_7;
  wire       [31:0]   addKernel_38_A_8;
  wire       [31:0]   addKernel_39_A_0;
  wire       [31:0]   addKernel_39_A_1;
  wire       [31:0]   addKernel_39_A_2;
  wire       [31:0]   addKernel_39_A_3;
  wire       [31:0]   addKernel_39_A_4;
  wire       [31:0]   addKernel_39_A_5;
  wire       [31:0]   addKernel_39_A_6;
  wire       [31:0]   addKernel_39_A_7;
  wire       [31:0]   addKernel_39_A_8;
  wire       [31:0]   addKernel_40_A_0;
  wire       [31:0]   addKernel_40_A_1;
  wire       [31:0]   addKernel_40_A_2;
  wire       [31:0]   addKernel_40_A_3;
  wire       [31:0]   addKernel_40_A_4;
  wire       [31:0]   addKernel_40_A_5;
  wire       [31:0]   addKernel_40_A_6;
  wire       [31:0]   addKernel_40_A_7;
  wire       [31:0]   addKernel_40_A_8;
  wire       [31:0]   addKernel_41_A_0;
  wire       [31:0]   addKernel_41_A_1;
  wire       [31:0]   addKernel_41_A_2;
  wire       [31:0]   addKernel_41_A_3;
  wire       [31:0]   addKernel_41_A_4;
  wire       [31:0]   addKernel_41_A_5;
  wire       [31:0]   addKernel_41_A_6;
  wire       [31:0]   addKernel_41_A_7;
  wire       [31:0]   addKernel_41_A_8;
  wire       [31:0]   addKernel_42_A_0;
  wire       [31:0]   addKernel_42_A_1;
  wire       [31:0]   addKernel_42_A_2;
  wire       [31:0]   addKernel_42_A_3;
  wire       [31:0]   addKernel_42_A_4;
  wire       [31:0]   addKernel_42_A_5;
  wire       [31:0]   addKernel_42_A_6;
  wire       [31:0]   addKernel_42_A_7;
  wire       [31:0]   addKernel_42_A_8;
  wire       [31:0]   addKernel_43_A_0;
  wire       [31:0]   addKernel_43_A_1;
  wire       [31:0]   addKernel_43_A_2;
  wire       [31:0]   addKernel_43_A_3;
  wire       [31:0]   addKernel_43_A_4;
  wire       [31:0]   addKernel_43_A_5;
  wire       [31:0]   addKernel_43_A_6;
  wire       [31:0]   addKernel_43_A_7;
  wire       [31:0]   addKernel_43_A_8;
  wire       [31:0]   addKernel_44_A_0;
  wire       [31:0]   addKernel_44_A_1;
  wire       [31:0]   addKernel_44_A_2;
  wire       [31:0]   addKernel_44_A_3;
  wire       [31:0]   addKernel_44_A_4;
  wire       [31:0]   addKernel_44_A_5;
  wire       [31:0]   addKernel_44_A_6;
  wire       [31:0]   addKernel_44_A_7;
  wire       [31:0]   addKernel_44_A_8;
  wire       [31:0]   addKernel_45_A_0;
  wire       [31:0]   addKernel_45_A_1;
  wire       [31:0]   addKernel_45_A_2;
  wire       [31:0]   addKernel_45_A_3;
  wire       [31:0]   addKernel_45_A_4;
  wire       [31:0]   addKernel_45_A_5;
  wire       [31:0]   addKernel_45_A_6;
  wire       [31:0]   addKernel_45_A_7;
  wire       [31:0]   addKernel_45_A_8;
  wire       [31:0]   addKernel_46_A_0;
  wire       [31:0]   addKernel_46_A_1;
  wire       [31:0]   addKernel_46_A_2;
  wire       [31:0]   addKernel_46_A_3;
  wire       [31:0]   addKernel_46_A_4;
  wire       [31:0]   addKernel_46_A_5;
  wire       [31:0]   addKernel_46_A_6;
  wire       [31:0]   addKernel_46_A_7;
  wire       [31:0]   addKernel_46_A_8;
  wire       [31:0]   addKernel_47_A_0;
  wire       [31:0]   addKernel_47_A_1;
  wire       [31:0]   addKernel_47_A_2;
  wire       [31:0]   addKernel_47_A_3;
  wire       [31:0]   addKernel_47_A_4;
  wire       [31:0]   addKernel_47_A_5;
  wire       [31:0]   addKernel_47_A_6;
  wire       [31:0]   addKernel_47_A_7;
  wire       [31:0]   addKernel_47_A_8;
  wire       [31:0]   addKernel_48_A_0;
  wire       [31:0]   addKernel_48_A_1;
  wire       [31:0]   addKernel_48_A_2;
  wire       [31:0]   addKernel_48_A_3;
  wire       [31:0]   addKernel_48_A_4;
  wire       [31:0]   addKernel_48_A_5;
  wire       [31:0]   addKernel_48_A_6;
  wire       [31:0]   addKernel_48_A_7;
  wire       [31:0]   addKernel_48_A_8;
  wire       [31:0]   addKernel_49_A_0;
  wire       [31:0]   addKernel_49_A_1;
  wire       [31:0]   addKernel_49_A_2;
  wire       [31:0]   addKernel_49_A_3;
  wire       [31:0]   addKernel_49_A_4;
  wire       [31:0]   addKernel_49_A_5;
  wire       [31:0]   addKernel_49_A_6;
  wire       [31:0]   addKernel_49_A_7;
  wire       [31:0]   addKernel_49_A_8;
  wire       [31:0]   addKernel_50_A_0;
  wire       [31:0]   addKernel_50_A_1;
  wire       [31:0]   addKernel_50_A_2;
  wire       [31:0]   addKernel_50_A_3;
  wire       [31:0]   addKernel_50_A_4;
  wire       [31:0]   addKernel_50_A_5;
  wire       [31:0]   addKernel_50_A_6;
  wire       [31:0]   addKernel_50_A_7;
  wire       [31:0]   addKernel_50_A_8;
  wire       [31:0]   addKernel_51_A_0;
  wire       [31:0]   addKernel_51_A_1;
  wire       [31:0]   addKernel_51_A_2;
  wire       [31:0]   addKernel_51_A_3;
  wire       [31:0]   addKernel_51_A_4;
  wire       [31:0]   addKernel_51_A_5;
  wire       [31:0]   addKernel_51_A_6;
  wire       [31:0]   addKernel_51_A_7;
  wire       [31:0]   addKernel_51_A_8;
  wire       [31:0]   addKernel_52_A_0;
  wire       [31:0]   addKernel_52_A_1;
  wire       [31:0]   addKernel_52_A_2;
  wire       [31:0]   addKernel_52_A_3;
  wire       [31:0]   addKernel_52_A_4;
  wire       [31:0]   addKernel_52_A_5;
  wire       [31:0]   addKernel_52_A_6;
  wire       [31:0]   addKernel_52_A_7;
  wire       [31:0]   addKernel_52_A_8;
  wire       [31:0]   addKernel_53_A_0;
  wire       [31:0]   addKernel_53_A_1;
  wire       [31:0]   addKernel_53_A_2;
  wire       [31:0]   addKernel_53_A_3;
  wire       [31:0]   addKernel_53_A_4;
  wire       [31:0]   addKernel_53_A_5;
  wire       [31:0]   addKernel_53_A_6;
  wire       [31:0]   addKernel_53_A_7;
  wire       [31:0]   addKernel_53_A_8;
  wire       [31:0]   addKernel_54_A_0;
  wire       [31:0]   addKernel_54_A_1;
  wire       [31:0]   addKernel_54_A_2;
  wire       [31:0]   addKernel_54_A_3;
  wire       [31:0]   addKernel_54_A_4;
  wire       [31:0]   addKernel_54_A_5;
  wire       [31:0]   addKernel_54_A_6;
  wire       [31:0]   addKernel_54_A_7;
  wire       [31:0]   addKernel_54_A_8;
  wire       [31:0]   addKernel_55_A_0;
  wire       [31:0]   addKernel_55_A_1;
  wire       [31:0]   addKernel_55_A_2;
  wire       [31:0]   addKernel_55_A_3;
  wire       [31:0]   addKernel_55_A_4;
  wire       [31:0]   addKernel_55_A_5;
  wire       [31:0]   addKernel_55_A_6;
  wire       [31:0]   addKernel_55_A_7;
  wire       [31:0]   addKernel_55_A_8;
  wire       [31:0]   addKernel_56_A_0;
  wire       [31:0]   addKernel_56_A_1;
  wire       [31:0]   addKernel_56_A_2;
  wire       [31:0]   addKernel_56_A_3;
  wire       [31:0]   addKernel_56_A_4;
  wire       [31:0]   addKernel_56_A_5;
  wire       [31:0]   addKernel_56_A_6;
  wire       [31:0]   addKernel_56_A_7;
  wire       [31:0]   addKernel_56_A_8;
  wire       [31:0]   addKernel_57_A_0;
  wire       [31:0]   addKernel_57_A_1;
  wire       [31:0]   addKernel_57_A_2;
  wire       [31:0]   addKernel_57_A_3;
  wire       [31:0]   addKernel_57_A_4;
  wire       [31:0]   addKernel_57_A_5;
  wire       [31:0]   addKernel_57_A_6;
  wire       [31:0]   addKernel_57_A_7;
  wire       [31:0]   addKernel_57_A_8;
  wire       [31:0]   addKernel_58_A_0;
  wire       [31:0]   addKernel_58_A_1;
  wire       [31:0]   addKernel_58_A_2;
  wire       [31:0]   addKernel_58_A_3;
  wire       [31:0]   addKernel_58_A_4;
  wire       [31:0]   addKernel_58_A_5;
  wire       [31:0]   addKernel_58_A_6;
  wire       [31:0]   addKernel_58_A_7;
  wire       [31:0]   addKernel_58_A_8;
  wire       [31:0]   addKernel_59_A_0;
  wire       [31:0]   addKernel_59_A_1;
  wire       [31:0]   addKernel_59_A_2;
  wire       [31:0]   addKernel_59_A_3;
  wire       [31:0]   addKernel_59_A_4;
  wire       [31:0]   addKernel_59_A_5;
  wire       [31:0]   addKernel_59_A_6;
  wire       [31:0]   addKernel_59_A_7;
  wire       [31:0]   addKernel_59_A_8;
  wire       [31:0]   addKernel_60_A_0;
  wire       [31:0]   addKernel_60_A_1;
  wire       [31:0]   addKernel_60_A_2;
  wire       [31:0]   addKernel_60_A_3;
  wire       [31:0]   addKernel_60_A_4;
  wire       [31:0]   addKernel_60_A_5;
  wire       [31:0]   addKernel_60_A_6;
  wire       [31:0]   addKernel_60_A_7;
  wire       [31:0]   addKernel_60_A_8;
  wire       [31:0]   addKernel_61_A_0;
  wire       [31:0]   addKernel_61_A_1;
  wire       [31:0]   addKernel_61_A_2;
  wire       [31:0]   addKernel_61_A_3;
  wire       [31:0]   addKernel_61_A_4;
  wire       [31:0]   addKernel_61_A_5;
  wire       [31:0]   addKernel_61_A_6;
  wire       [31:0]   addKernel_61_A_7;
  wire       [31:0]   addKernel_61_A_8;
  wire       [31:0]   addKernel_62_A_0;
  wire       [31:0]   addKernel_62_A_1;
  wire       [31:0]   addKernel_62_A_2;
  wire       [31:0]   addKernel_62_A_3;
  wire       [31:0]   addKernel_62_A_4;
  wire       [31:0]   addKernel_62_A_5;
  wire       [31:0]   addKernel_62_A_6;
  wire       [31:0]   addKernel_62_A_7;
  wire       [31:0]   addKernel_62_A_8;
  wire       [31:0]   addKernel_63_A_0;
  wire       [31:0]   addKernel_63_A_1;
  wire       [31:0]   addKernel_63_A_2;
  wire       [31:0]   addKernel_63_A_3;
  wire       [31:0]   addKernel_63_A_4;
  wire       [31:0]   addKernel_63_A_5;
  wire       [31:0]   addKernel_63_A_6;
  wire       [31:0]   addKernel_63_A_7;
  wire       [31:0]   addKernel_63_A_8;
  wire       [31:0]   addKernel_64_A_0;
  wire       [31:0]   addKernel_64_A_1;
  wire       [31:0]   addKernel_64_A_2;
  wire       [31:0]   addKernel_64_A_3;
  wire       [31:0]   addKernel_64_A_4;
  wire       [31:0]   addKernel_64_A_5;
  wire       [31:0]   addKernel_64_A_6;
  wire       [31:0]   addKernel_64_A_7;
  wire       [31:0]   addKernel_64_A_8;
  wire       [31:0]   addKernel_65_A_0;
  wire       [31:0]   addKernel_65_A_1;
  wire       [31:0]   addKernel_65_A_2;
  wire       [31:0]   addKernel_65_A_3;
  wire       [31:0]   addKernel_65_A_4;
  wire       [31:0]   addKernel_65_A_5;
  wire       [31:0]   addKernel_65_A_6;
  wire       [31:0]   addKernel_65_A_7;
  wire       [31:0]   addKernel_65_A_8;
  wire       [31:0]   addKernel_66_A_0;
  wire       [31:0]   addKernel_66_A_1;
  wire       [31:0]   addKernel_66_A_2;
  wire       [31:0]   addKernel_66_A_3;
  wire       [31:0]   addKernel_66_A_4;
  wire       [31:0]   addKernel_66_A_5;
  wire       [31:0]   addKernel_66_A_6;
  wire       [31:0]   addKernel_66_A_7;
  wire       [31:0]   addKernel_66_A_8;
  wire       [31:0]   addKernel_67_A_0;
  wire       [31:0]   addKernel_67_A_1;
  wire       [31:0]   addKernel_67_A_2;
  wire       [31:0]   addKernel_67_A_3;
  wire       [31:0]   addKernel_67_A_4;
  wire       [31:0]   addKernel_67_A_5;
  wire       [31:0]   addKernel_67_A_6;
  wire       [31:0]   addKernel_67_A_7;
  wire       [31:0]   addKernel_67_A_8;
  wire       [31:0]   addKernel_68_A_0;
  wire       [31:0]   addKernel_68_A_1;
  wire       [31:0]   addKernel_68_A_2;
  wire       [31:0]   addKernel_68_A_3;
  wire       [31:0]   addKernel_68_A_4;
  wire       [31:0]   addKernel_68_A_5;
  wire       [31:0]   addKernel_68_A_6;
  wire       [31:0]   addKernel_68_A_7;
  wire       [31:0]   addKernel_68_A_8;
  wire       [31:0]   addKernel_69_A_0;
  wire       [31:0]   addKernel_69_A_1;
  wire       [31:0]   addKernel_69_A_2;
  wire       [31:0]   addKernel_69_A_3;
  wire       [31:0]   addKernel_69_A_4;
  wire       [31:0]   addKernel_69_A_5;
  wire       [31:0]   addKernel_69_A_6;
  wire       [31:0]   addKernel_69_A_7;
  wire       [31:0]   addKernel_69_A_8;
  wire       [31:0]   addKernel_70_A_0;
  wire       [31:0]   addKernel_70_A_1;
  wire       [31:0]   addKernel_70_A_2;
  wire       [31:0]   addKernel_70_A_3;
  wire       [31:0]   addKernel_70_A_4;
  wire       [31:0]   addKernel_70_A_5;
  wire       [31:0]   addKernel_70_A_6;
  wire       [31:0]   addKernel_70_A_7;
  wire       [31:0]   addKernel_70_A_8;
  wire       [31:0]   addKernel_71_A_0;
  wire       [31:0]   addKernel_71_A_1;
  wire       [31:0]   addKernel_71_A_2;
  wire       [31:0]   addKernel_71_A_3;
  wire       [31:0]   addKernel_71_A_4;
  wire       [31:0]   addKernel_71_A_5;
  wire       [31:0]   addKernel_71_A_6;
  wire       [31:0]   addKernel_71_A_7;
  wire       [31:0]   addKernel_71_A_8;
  wire       [31:0]   addKernel_72_A_0;
  wire       [31:0]   addKernel_72_A_1;
  wire       [31:0]   addKernel_72_A_2;
  wire       [31:0]   addKernel_72_A_3;
  wire       [31:0]   addKernel_72_A_4;
  wire       [31:0]   addKernel_72_A_5;
  wire       [31:0]   addKernel_72_A_6;
  wire       [31:0]   addKernel_72_A_7;
  wire       [31:0]   addKernel_72_A_8;
  wire       [31:0]   addKernel_73_A_0;
  wire       [31:0]   addKernel_73_A_1;
  wire       [31:0]   addKernel_73_A_2;
  wire       [31:0]   addKernel_73_A_3;
  wire       [31:0]   addKernel_73_A_4;
  wire       [31:0]   addKernel_73_A_5;
  wire       [31:0]   addKernel_73_A_6;
  wire       [31:0]   addKernel_73_A_7;
  wire       [31:0]   addKernel_73_A_8;
  wire       [31:0]   addKernel_74_A_0;
  wire       [31:0]   addKernel_74_A_1;
  wire       [31:0]   addKernel_74_A_2;
  wire       [31:0]   addKernel_74_A_3;
  wire       [31:0]   addKernel_74_A_4;
  wire       [31:0]   addKernel_74_A_5;
  wire       [31:0]   addKernel_74_A_6;
  wire       [31:0]   addKernel_74_A_7;
  wire       [31:0]   addKernel_74_A_8;
  wire       [31:0]   addKernel_75_A_0;
  wire       [31:0]   addKernel_75_A_1;
  wire       [31:0]   addKernel_75_A_2;
  wire       [31:0]   addKernel_75_A_3;
  wire       [31:0]   addKernel_75_A_4;
  wire       [31:0]   addKernel_75_A_5;
  wire       [31:0]   addKernel_75_A_6;
  wire       [31:0]   addKernel_75_A_7;
  wire       [31:0]   addKernel_75_A_8;
  wire       [31:0]   addKernel_76_A_0;
  wire       [31:0]   addKernel_76_A_1;
  wire       [31:0]   addKernel_76_A_2;
  wire       [31:0]   addKernel_76_A_3;
  wire       [31:0]   addKernel_76_A_4;
  wire       [31:0]   addKernel_76_A_5;
  wire       [31:0]   addKernel_76_A_6;
  wire       [31:0]   addKernel_76_A_7;
  wire       [31:0]   addKernel_76_A_8;
  wire       [31:0]   addKernel_77_A_0;
  wire       [31:0]   addKernel_77_A_1;
  wire       [31:0]   addKernel_77_A_2;
  wire       [31:0]   addKernel_77_A_3;
  wire       [31:0]   addKernel_77_A_4;
  wire       [31:0]   addKernel_77_A_5;
  wire       [31:0]   addKernel_77_A_6;
  wire       [31:0]   addKernel_77_A_7;
  wire       [31:0]   addKernel_77_A_8;
  wire       [31:0]   addKernel_78_A_0;
  wire       [31:0]   addKernel_78_A_1;
  wire       [31:0]   addKernel_78_A_2;
  wire       [31:0]   addKernel_78_A_3;
  wire       [31:0]   addKernel_78_A_4;
  wire       [31:0]   addKernel_78_A_5;
  wire       [31:0]   addKernel_78_A_6;
  wire       [31:0]   addKernel_78_A_7;
  wire       [31:0]   addKernel_78_A_8;
  wire       [31:0]   addKernel_79_A_0;
  wire       [31:0]   addKernel_79_A_1;
  wire       [31:0]   addKernel_79_A_2;
  wire       [31:0]   addKernel_79_A_3;
  wire       [31:0]   addKernel_79_A_4;
  wire       [31:0]   addKernel_79_A_5;
  wire       [31:0]   addKernel_79_A_6;
  wire       [31:0]   addKernel_79_A_7;
  wire       [31:0]   addKernel_79_A_8;
  wire       [31:0]   addKernel_80_A_0;
  wire       [31:0]   addKernel_80_A_1;
  wire       [31:0]   addKernel_80_A_2;
  wire       [31:0]   addKernel_80_A_3;
  wire       [31:0]   addKernel_80_A_4;
  wire       [31:0]   addKernel_80_A_5;
  wire       [31:0]   addKernel_80_A_6;
  wire       [31:0]   addKernel_80_A_7;
  wire       [31:0]   addKernel_80_A_8;
  wire       [31:0]   addKernel_81_A_0;
  wire       [31:0]   addKernel_81_A_1;
  wire       [31:0]   addKernel_81_A_2;
  wire       [31:0]   addKernel_81_A_3;
  wire       [31:0]   addKernel_81_A_4;
  wire       [31:0]   addKernel_81_A_5;
  wire       [31:0]   addKernel_81_A_6;
  wire       [31:0]   addKernel_81_A_7;
  wire       [31:0]   addKernel_81_A_8;
  wire       [31:0]   addKernel_82_A_0;
  wire       [31:0]   addKernel_82_A_1;
  wire       [31:0]   addKernel_82_A_2;
  wire       [31:0]   addKernel_82_A_3;
  wire       [31:0]   addKernel_82_A_4;
  wire       [31:0]   addKernel_82_A_5;
  wire       [31:0]   addKernel_82_A_6;
  wire       [31:0]   addKernel_82_A_7;
  wire       [31:0]   addKernel_82_A_8;
  wire       [31:0]   addKernel_83_A_0;
  wire       [31:0]   addKernel_83_A_1;
  wire       [31:0]   addKernel_83_A_2;
  wire       [31:0]   addKernel_83_A_3;
  wire       [31:0]   addKernel_83_A_4;
  wire       [31:0]   addKernel_83_A_5;
  wire       [31:0]   addKernel_83_A_6;
  wire       [31:0]   addKernel_83_A_7;
  wire       [31:0]   addKernel_83_A_8;
  wire       [31:0]   addKernel_84_A_0;
  wire       [31:0]   addKernel_84_A_1;
  wire       [31:0]   addKernel_84_A_2;
  wire       [31:0]   addKernel_84_A_3;
  wire       [31:0]   addKernel_84_A_4;
  wire       [31:0]   addKernel_84_A_5;
  wire       [31:0]   addKernel_84_A_6;
  wire       [31:0]   addKernel_84_A_7;
  wire       [31:0]   addKernel_84_A_8;
  wire       [31:0]   addKernel_85_A_0;
  wire       [31:0]   addKernel_85_A_1;
  wire       [31:0]   addKernel_85_A_2;
  wire       [31:0]   addKernel_85_A_3;
  wire       [31:0]   addKernel_85_A_4;
  wire       [31:0]   addKernel_85_A_5;
  wire       [31:0]   addKernel_85_A_6;
  wire       [31:0]   addKernel_85_A_7;
  wire       [31:0]   addKernel_85_A_8;
  wire       [31:0]   addKernel_86_A_0;
  wire       [31:0]   addKernel_86_A_1;
  wire       [31:0]   addKernel_86_A_2;
  wire       [31:0]   addKernel_86_A_3;
  wire       [31:0]   addKernel_86_A_4;
  wire       [31:0]   addKernel_86_A_5;
  wire       [31:0]   addKernel_86_A_6;
  wire       [31:0]   addKernel_86_A_7;
  wire       [31:0]   addKernel_86_A_8;
  wire       [31:0]   addKernel_87_A_0;
  wire       [31:0]   addKernel_87_A_1;
  wire       [31:0]   addKernel_87_A_2;
  wire       [31:0]   addKernel_87_A_3;
  wire       [31:0]   addKernel_87_A_4;
  wire       [31:0]   addKernel_87_A_5;
  wire       [31:0]   addKernel_87_A_6;
  wire       [31:0]   addKernel_87_A_7;
  wire       [31:0]   addKernel_87_A_8;
  wire       [31:0]   addKernel_88_A_0;
  wire       [31:0]   addKernel_88_A_1;
  wire       [31:0]   addKernel_88_A_2;
  wire       [31:0]   addKernel_88_A_3;
  wire       [31:0]   addKernel_88_A_4;
  wire       [31:0]   addKernel_88_A_5;
  wire       [31:0]   addKernel_88_A_6;
  wire       [31:0]   addKernel_88_A_7;
  wire       [31:0]   addKernel_88_A_8;
  wire       [31:0]   addKernel_89_A_0;
  wire       [31:0]   addKernel_89_A_1;
  wire       [31:0]   addKernel_89_A_2;
  wire       [31:0]   addKernel_89_A_3;
  wire       [31:0]   addKernel_89_A_4;
  wire       [31:0]   addKernel_89_A_5;
  wire       [31:0]   addKernel_89_A_6;
  wire       [31:0]   addKernel_89_A_7;
  wire       [31:0]   addKernel_89_A_8;
  wire       [31:0]   addKernel_90_A_0;
  wire       [31:0]   addKernel_90_A_1;
  wire       [31:0]   addKernel_90_A_2;
  wire       [31:0]   addKernel_90_A_3;
  wire       [31:0]   addKernel_90_A_4;
  wire       [31:0]   addKernel_90_A_5;
  wire       [31:0]   addKernel_90_A_6;
  wire       [31:0]   addKernel_90_A_7;
  wire       [31:0]   addKernel_90_A_8;
  wire       [31:0]   addKernel_91_A_0;
  wire       [31:0]   addKernel_91_A_1;
  wire       [31:0]   addKernel_91_A_2;
  wire       [31:0]   addKernel_91_A_3;
  wire       [31:0]   addKernel_91_A_4;
  wire       [31:0]   addKernel_91_A_5;
  wire       [31:0]   addKernel_91_A_6;
  wire       [31:0]   addKernel_91_A_7;
  wire       [31:0]   addKernel_91_A_8;
  wire       [31:0]   addKernel_92_A_0;
  wire       [31:0]   addKernel_92_A_1;
  wire       [31:0]   addKernel_92_A_2;
  wire       [31:0]   addKernel_92_A_3;
  wire       [31:0]   addKernel_92_A_4;
  wire       [31:0]   addKernel_92_A_5;
  wire       [31:0]   addKernel_92_A_6;
  wire       [31:0]   addKernel_92_A_7;
  wire       [31:0]   addKernel_92_A_8;
  wire       [31:0]   addKernel_93_A_0;
  wire       [31:0]   addKernel_93_A_1;
  wire       [31:0]   addKernel_93_A_2;
  wire       [31:0]   addKernel_93_A_3;
  wire       [31:0]   addKernel_93_A_4;
  wire       [31:0]   addKernel_93_A_5;
  wire       [31:0]   addKernel_93_A_6;
  wire       [31:0]   addKernel_93_A_7;
  wire       [31:0]   addKernel_93_A_8;
  wire       [31:0]   addKernel_94_A_0;
  wire       [31:0]   addKernel_94_A_1;
  wire       [31:0]   addKernel_94_A_2;
  wire       [31:0]   addKernel_94_A_3;
  wire       [31:0]   addKernel_94_A_4;
  wire       [31:0]   addKernel_94_A_5;
  wire       [31:0]   addKernel_94_A_6;
  wire       [31:0]   addKernel_94_A_7;
  wire       [31:0]   addKernel_94_A_8;
  wire       [31:0]   addKernel_95_A_0;
  wire       [31:0]   addKernel_95_A_1;
  wire       [31:0]   addKernel_95_A_2;
  wire       [31:0]   addKernel_95_A_3;
  wire       [31:0]   addKernel_95_A_4;
  wire       [31:0]   addKernel_95_A_5;
  wire       [31:0]   addKernel_95_A_6;
  wire       [31:0]   addKernel_95_A_7;
  wire       [31:0]   addKernel_95_A_8;
  wire       [31:0]   addKernel_96_A_0;
  wire       [31:0]   addKernel_96_A_1;
  wire       [31:0]   addKernel_96_A_2;
  wire       [31:0]   addKernel_96_A_3;
  wire       [31:0]   addKernel_96_A_4;
  wire       [31:0]   addKernel_96_A_5;
  wire       [31:0]   addKernel_96_A_6;
  wire       [31:0]   addKernel_96_A_7;
  wire       [31:0]   addKernel_96_A_8;
  wire       [31:0]   addKernel_97_A_0;
  wire       [31:0]   addKernel_97_A_1;
  wire       [31:0]   addKernel_97_A_2;
  wire       [31:0]   addKernel_97_A_3;
  wire       [31:0]   addKernel_97_A_4;
  wire       [31:0]   addKernel_97_A_5;
  wire       [31:0]   addKernel_97_A_6;
  wire       [31:0]   addKernel_97_A_7;
  wire       [31:0]   addKernel_97_A_8;
  wire       [31:0]   addKernel_98_A_0;
  wire       [31:0]   addKernel_98_A_1;
  wire       [31:0]   addKernel_98_A_2;
  wire       [31:0]   addKernel_98_A_3;
  wire       [31:0]   addKernel_98_A_4;
  wire       [31:0]   addKernel_98_A_5;
  wire       [31:0]   addKernel_98_A_6;
  wire       [31:0]   addKernel_98_A_7;
  wire       [31:0]   addKernel_98_A_8;
  wire       [31:0]   addKernel_99_A_0;
  wire       [31:0]   addKernel_99_A_1;
  wire       [31:0]   addKernel_99_A_2;
  wire       [31:0]   addKernel_99_A_3;
  wire       [31:0]   addKernel_99_A_4;
  wire       [31:0]   addKernel_99_A_5;
  wire       [31:0]   addKernel_99_A_6;
  wire       [31:0]   addKernel_99_A_7;
  wire       [31:0]   addKernel_99_A_8;
  wire       [31:0]   addKernel_100_A_0;
  wire       [31:0]   addKernel_100_A_1;
  wire       [31:0]   addKernel_100_A_2;
  wire       [31:0]   addKernel_100_A_3;
  wire       [31:0]   addKernel_100_A_4;
  wire       [31:0]   addKernel_100_A_5;
  wire       [31:0]   addKernel_100_A_6;
  wire       [31:0]   addKernel_100_A_7;
  wire       [31:0]   addKernel_100_A_8;
  wire       [31:0]   addKernel_101_A_0;
  wire       [31:0]   addKernel_101_A_1;
  wire       [31:0]   addKernel_101_A_2;
  wire       [31:0]   addKernel_101_A_3;
  wire       [31:0]   addKernel_101_A_4;
  wire       [31:0]   addKernel_101_A_5;
  wire       [31:0]   addKernel_101_A_6;
  wire       [31:0]   addKernel_101_A_7;
  wire       [31:0]   addKernel_101_A_8;
  wire       [31:0]   addKernel_102_A_0;
  wire       [31:0]   addKernel_102_A_1;
  wire       [31:0]   addKernel_102_A_2;
  wire       [31:0]   addKernel_102_A_3;
  wire       [31:0]   addKernel_102_A_4;
  wire       [31:0]   addKernel_102_A_5;
  wire       [31:0]   addKernel_102_A_6;
  wire       [31:0]   addKernel_102_A_7;
  wire       [31:0]   addKernel_102_A_8;
  wire       [31:0]   addKernel_103_A_0;
  wire       [31:0]   addKernel_103_A_1;
  wire       [31:0]   addKernel_103_A_2;
  wire       [31:0]   addKernel_103_A_3;
  wire       [31:0]   addKernel_103_A_4;
  wire       [31:0]   addKernel_103_A_5;
  wire       [31:0]   addKernel_103_A_6;
  wire       [31:0]   addKernel_103_A_7;
  wire       [31:0]   addKernel_103_A_8;
  wire       [31:0]   addKernel_104_A_0;
  wire       [31:0]   addKernel_104_A_1;
  wire       [31:0]   addKernel_104_A_2;
  wire       [31:0]   addKernel_104_A_3;
  wire       [31:0]   addKernel_104_A_4;
  wire       [31:0]   addKernel_104_A_5;
  wire       [31:0]   addKernel_104_A_6;
  wire       [31:0]   addKernel_104_A_7;
  wire       [31:0]   addKernel_104_A_8;
  wire       [31:0]   addKernel_105_A_0;
  wire       [31:0]   addKernel_105_A_1;
  wire       [31:0]   addKernel_105_A_2;
  wire       [31:0]   addKernel_105_A_3;
  wire       [31:0]   addKernel_105_A_4;
  wire       [31:0]   addKernel_105_A_5;
  wire       [31:0]   addKernel_105_A_6;
  wire       [31:0]   addKernel_105_A_7;
  wire       [31:0]   addKernel_105_A_8;
  wire       [31:0]   addKernel_106_A_0;
  wire       [31:0]   addKernel_106_A_1;
  wire       [31:0]   addKernel_106_A_2;
  wire       [31:0]   addKernel_106_A_3;
  wire       [31:0]   addKernel_106_A_4;
  wire       [31:0]   addKernel_106_A_5;
  wire       [31:0]   addKernel_106_A_6;
  wire       [31:0]   addKernel_106_A_7;
  wire       [31:0]   addKernel_106_A_8;
  wire       [31:0]   addKernel_107_A_0;
  wire       [31:0]   addKernel_107_A_1;
  wire       [31:0]   addKernel_107_A_2;
  wire       [31:0]   addKernel_107_A_3;
  wire       [31:0]   addKernel_107_A_4;
  wire       [31:0]   addKernel_107_A_5;
  wire       [31:0]   addKernel_107_A_6;
  wire       [31:0]   addKernel_107_A_7;
  wire       [31:0]   addKernel_107_A_8;
  wire       [31:0]   addKernel_108_A_0;
  wire       [31:0]   addKernel_108_A_1;
  wire       [31:0]   addKernel_108_A_2;
  wire       [31:0]   addKernel_108_A_3;
  wire       [31:0]   addKernel_108_A_4;
  wire       [31:0]   addKernel_108_A_5;
  wire       [31:0]   addKernel_108_A_6;
  wire       [31:0]   addKernel_108_A_7;
  wire       [31:0]   addKernel_108_A_8;
  wire       [31:0]   addKernel_109_A_0;
  wire       [31:0]   addKernel_109_A_1;
  wire       [31:0]   addKernel_109_A_2;
  wire       [31:0]   addKernel_109_A_3;
  wire       [31:0]   addKernel_109_A_4;
  wire       [31:0]   addKernel_109_A_5;
  wire       [31:0]   addKernel_109_A_6;
  wire       [31:0]   addKernel_109_A_7;
  wire       [31:0]   addKernel_109_A_8;
  wire       [31:0]   addKernel_110_A_0;
  wire       [31:0]   addKernel_110_A_1;
  wire       [31:0]   addKernel_110_A_2;
  wire       [31:0]   addKernel_110_A_3;
  wire       [31:0]   addKernel_110_A_4;
  wire       [31:0]   addKernel_110_A_5;
  wire       [31:0]   addKernel_110_A_6;
  wire       [31:0]   addKernel_110_A_7;
  wire       [31:0]   addKernel_110_A_8;
  wire       [31:0]   addKernel_111_A_0;
  wire       [31:0]   addKernel_111_A_1;
  wire       [31:0]   addKernel_111_A_2;
  wire       [31:0]   addKernel_111_A_3;
  wire       [31:0]   addKernel_111_A_4;
  wire       [31:0]   addKernel_111_A_5;
  wire       [31:0]   addKernel_111_A_6;
  wire       [31:0]   addKernel_111_A_7;
  wire       [31:0]   addKernel_111_A_8;
  wire       [31:0]   addKernel_112_A_0;
  wire       [31:0]   addKernel_112_A_1;
  wire       [31:0]   addKernel_112_A_2;
  wire       [31:0]   addKernel_112_A_3;
  wire       [31:0]   addKernel_112_A_4;
  wire       [31:0]   addKernel_112_A_5;
  wire       [31:0]   addKernel_112_A_6;
  wire       [31:0]   addKernel_112_A_7;
  wire       [31:0]   addKernel_112_A_8;
  wire       [31:0]   addKernel_113_A_0;
  wire       [31:0]   addKernel_113_A_1;
  wire       [31:0]   addKernel_113_A_2;
  wire       [31:0]   addKernel_113_A_3;
  wire       [31:0]   addKernel_113_A_4;
  wire       [31:0]   addKernel_113_A_5;
  wire       [31:0]   addKernel_113_A_6;
  wire       [31:0]   addKernel_113_A_7;
  wire       [31:0]   addKernel_113_A_8;
  wire       [31:0]   addKernel_114_A_0;
  wire       [31:0]   addKernel_114_A_1;
  wire       [31:0]   addKernel_114_A_2;
  wire       [31:0]   addKernel_114_A_3;
  wire       [31:0]   addKernel_114_A_4;
  wire       [31:0]   addKernel_114_A_5;
  wire       [31:0]   addKernel_114_A_6;
  wire       [31:0]   addKernel_114_A_7;
  wire       [31:0]   addKernel_114_A_8;
  wire       [31:0]   addKernel_115_A_0;
  wire       [31:0]   addKernel_115_A_1;
  wire       [31:0]   addKernel_115_A_2;
  wire       [31:0]   addKernel_115_A_3;
  wire       [31:0]   addKernel_115_A_4;
  wire       [31:0]   addKernel_115_A_5;
  wire       [31:0]   addKernel_115_A_6;
  wire       [31:0]   addKernel_115_A_7;
  wire       [31:0]   addKernel_115_A_8;
  wire       [31:0]   addKernel_116_A_0;
  wire       [31:0]   addKernel_116_A_1;
  wire       [31:0]   addKernel_116_A_2;
  wire       [31:0]   addKernel_116_A_3;
  wire       [31:0]   addKernel_116_A_4;
  wire       [31:0]   addKernel_116_A_5;
  wire       [31:0]   addKernel_116_A_6;
  wire       [31:0]   addKernel_116_A_7;
  wire       [31:0]   addKernel_116_A_8;
  wire       [31:0]   addKernel_117_A_0;
  wire       [31:0]   addKernel_117_A_1;
  wire       [31:0]   addKernel_117_A_2;
  wire       [31:0]   addKernel_117_A_3;
  wire       [31:0]   addKernel_117_A_4;
  wire       [31:0]   addKernel_117_A_5;
  wire       [31:0]   addKernel_117_A_6;
  wire       [31:0]   addKernel_117_A_7;
  wire       [31:0]   addKernel_117_A_8;
  wire       [31:0]   addKernel_118_A_0;
  wire       [31:0]   addKernel_118_A_1;
  wire       [31:0]   addKernel_118_A_2;
  wire       [31:0]   addKernel_118_A_3;
  wire       [31:0]   addKernel_118_A_4;
  wire       [31:0]   addKernel_118_A_5;
  wire       [31:0]   addKernel_118_A_6;
  wire       [31:0]   addKernel_118_A_7;
  wire       [31:0]   addKernel_118_A_8;
  wire       [31:0]   addKernel_119_A_0;
  wire       [31:0]   addKernel_119_A_1;
  wire       [31:0]   addKernel_119_A_2;
  wire       [31:0]   addKernel_119_A_3;
  wire       [31:0]   addKernel_119_A_4;
  wire       [31:0]   addKernel_119_A_5;
  wire       [31:0]   addKernel_119_A_6;
  wire       [31:0]   addKernel_119_A_7;
  wire       [31:0]   addKernel_119_A_8;
  wire       [31:0]   addKernel_120_A_0;
  wire       [31:0]   addKernel_120_A_1;
  wire       [31:0]   addKernel_120_A_2;
  wire       [31:0]   addKernel_120_A_3;
  wire       [31:0]   addKernel_120_A_4;
  wire       [31:0]   addKernel_120_A_5;
  wire       [31:0]   addKernel_120_A_6;
  wire       [31:0]   addKernel_120_A_7;
  wire       [31:0]   addKernel_120_A_8;
  wire       [31:0]   addKernel_121_A_0;
  wire       [31:0]   addKernel_121_A_1;
  wire       [31:0]   addKernel_121_A_2;
  wire       [31:0]   addKernel_121_A_3;
  wire       [31:0]   addKernel_121_A_4;
  wire       [31:0]   addKernel_121_A_5;
  wire       [31:0]   addKernel_121_A_6;
  wire       [31:0]   addKernel_121_A_7;
  wire       [31:0]   addKernel_121_A_8;
  wire       [31:0]   addKernel_122_A_0;
  wire       [31:0]   addKernel_122_A_1;
  wire       [31:0]   addKernel_122_A_2;
  wire       [31:0]   addKernel_122_A_3;
  wire       [31:0]   addKernel_122_A_4;
  wire       [31:0]   addKernel_122_A_5;
  wire       [31:0]   addKernel_122_A_6;
  wire       [31:0]   addKernel_122_A_7;
  wire       [31:0]   addKernel_122_A_8;
  wire       [31:0]   addKernel_123_A_0;
  wire       [31:0]   addKernel_123_A_1;
  wire       [31:0]   addKernel_123_A_2;
  wire       [31:0]   addKernel_123_A_3;
  wire       [31:0]   addKernel_123_A_4;
  wire       [31:0]   addKernel_123_A_5;
  wire       [31:0]   addKernel_123_A_6;
  wire       [31:0]   addKernel_123_A_7;
  wire       [31:0]   addKernel_123_A_8;
  wire       [31:0]   addKernel_124_A_0;
  wire       [31:0]   addKernel_124_A_1;
  wire       [31:0]   addKernel_124_A_2;
  wire       [31:0]   addKernel_124_A_3;
  wire       [31:0]   addKernel_124_A_4;
  wire       [31:0]   addKernel_124_A_5;
  wire       [31:0]   addKernel_124_A_6;
  wire       [31:0]   addKernel_124_A_7;
  wire       [31:0]   addKernel_124_A_8;
  wire       [31:0]   addKernel_125_A_0;
  wire       [31:0]   addKernel_125_A_1;
  wire       [31:0]   addKernel_125_A_2;
  wire       [31:0]   addKernel_125_A_3;
  wire       [31:0]   addKernel_125_A_4;
  wire       [31:0]   addKernel_125_A_5;
  wire       [31:0]   addKernel_125_A_6;
  wire       [31:0]   addKernel_125_A_7;
  wire       [31:0]   addKernel_125_A_8;
  wire       [31:0]   addKernel_126_A_0;
  wire       [31:0]   addKernel_126_A_1;
  wire       [31:0]   addKernel_126_A_2;
  wire       [31:0]   addKernel_126_A_3;
  wire       [31:0]   addKernel_126_A_4;
  wire       [31:0]   addKernel_126_A_5;
  wire       [31:0]   addKernel_126_A_6;
  wire       [31:0]   addKernel_126_A_7;
  wire       [31:0]   addKernel_126_A_8;
  wire       [31:0]   addKernel_127_A_0;
  wire       [31:0]   addKernel_127_A_1;
  wire       [31:0]   addKernel_127_A_2;
  wire       [31:0]   addKernel_127_A_3;
  wire       [31:0]   addKernel_127_A_4;
  wire       [31:0]   addKernel_127_A_5;
  wire       [31:0]   addKernel_127_A_6;
  wire       [31:0]   addKernel_127_A_7;
  wire       [31:0]   addKernel_127_A_8;
  wire       [23:0]   xAddChannelTimes_16_A;
  wire       [23:0]   xAddChannelTimes_17_A;
  wire       [23:0]   xAddChannelTimes_18_A;
  wire       [23:0]   xAddChannelTimes_19_A;
  wire       [23:0]   xAddChannelTimes_20_A;
  wire       [23:0]   xAddChannelTimes_21_A;
  wire       [23:0]   xAddChannelTimes_22_A;
  wire       [23:0]   xAddChannelTimes_23_A;
  wire       [23:0]   xAddChannelTimes_24_A;
  wire       [23:0]   xAddChannelTimes_25_A;
  wire       [23:0]   xAddChannelTimes_26_A;
  wire       [23:0]   xAddChannelTimes_27_A;
  wire       [23:0]   xAddChannelTimes_28_A;
  wire       [23:0]   xAddChannelTimes_29_A;
  wire       [23:0]   xAddChannelTimes_30_A;
  wire       [23:0]   xAddChannelTimes_31_A;
  reg        [127:0]  _zz__zz_1_port1;
  reg        [127:0]  _zz__zz_2_port1;
  reg        [127:0]  _zz__zz_3_port1;
  reg        [127:0]  _zz__zz_4_port1;
  reg        [127:0]  _zz__zz_5_port1;
  reg        [127:0]  _zz__zz_6_port1;
  reg        [127:0]  _zz__zz_7_port1;
  reg        [127:0]  _zz__zz_8_port1;
  reg        [127:0]  _zz__zz_9_port1;
  wire                channelIncr_1_sData_ready;
  wire                channelIncr_1_mData_valid;
  wire       [127:0]  channelIncr_1_mData_payload;
  wire                dataGenerate_1_sData_ready;
  wire                dataGenerate_1_mData_mData_0_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_0_payload;
  wire                dataGenerate_1_mData_mData_1_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_1_payload;
  wire                dataGenerate_1_mData_mData_2_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_2_payload;
  wire                dataGenerate_1_mData_mData_3_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_3_payload;
  wire                dataGenerate_1_mData_mData_4_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_4_payload;
  wire                dataGenerate_1_mData_mData_5_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_5_payload;
  wire                dataGenerate_1_mData_mData_6_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_6_payload;
  wire                dataGenerate_1_mData_mData_7_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_7_payload;
  wire                dataGenerate_1_mData_mData_8_valid;
  wire       [127:0]  dataGenerate_1_mData_mData_8_payload;
  wire                convComputeCtrl_1_mDataValid;
  wire                convComputeCtrl_1_normPreValid;
  wire       [4:0]    convComputeCtrl_1_featureMemReadAddr;
  wire       [4:0]    convComputeCtrl_1_featureMemWriteAddr;
  wire                convComputeCtrl_1_featureMemWriteReady;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_0;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_1;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_2;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_3;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_4;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_5;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_6;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_7;
  wire       [8:0]    convComputeCtrl_1_weightReadAddr_8;
  wire       [5:0]    convComputeCtrl_1_biasReadAddr;
  wire       [5:0]    convComputeCtrl_1_scaleReadAddr;
  wire       [5:0]    convComputeCtrl_1_shiftReadAddr;
  wire       [12:0]   convComputeCtrl_1_sCount;
  wire       [12:0]   convComputeCtrl_1_mCount;
  wire                loadWeight_1_sData_ready;
  wire       [2047:0] loadWeight_1_weightRead_0_data;
  wire       [2047:0] loadWeight_1_weightRead_1_data;
  wire       [2047:0] loadWeight_1_weightRead_2_data;
  wire       [2047:0] loadWeight_1_weightRead_3_data;
  wire       [2047:0] loadWeight_1_weightRead_4_data;
  wire       [2047:0] loadWeight_1_weightRead_5_data;
  wire       [2047:0] loadWeight_1_weightRead_6_data;
  wire       [2047:0] loadWeight_1_weightRead_7_data;
  wire       [2047:0] loadWeight_1_weightRead_8_data;
  wire       [511:0]  loadWeight_1_biasRead_data;
  wire       [511:0]  loadWeight_1_scaleRead_data;
  wire       [511:0]  loadWeight_1_shiftRead_data;
  wire                loadWeight_1_copyWeightDone;
  wire                waXpmSyncFifo_9_sReady;
  wire                waXpmSyncFifo_9_mReady;
  wire       [127:0]  waXpmSyncFifo_9_dout;
  wire       [127:0]  waXpmSyncFifo_10_dout;
  wire       [127:0]  waXpmSyncFifo_11_dout;
  wire       [127:0]  waXpmSyncFifo_12_dout;
  wire       [127:0]  waXpmSyncFifo_13_dout;
  wire       [127:0]  waXpmSyncFifo_14_dout;
  wire       [127:0]  waXpmSyncFifo_15_dout;
  wire       [127:0]  waXpmSyncFifo_16_dout;
  wire       [127:0]  waXpmSyncFifo_17_dout;
  wire       [31:0]   dSP_1_p;
  wire       [31:0]   dSP_2_p;
  wire       [31:0]   dSP_3_p;
  wire       [31:0]   dSP_4_p;
  wire       [31:0]   dSP_5_p;
  wire       [31:0]   dSP_6_p;
  wire       [31:0]   dSP_7_p;
  wire       [31:0]   dSP_8_p;
  wire       [31:0]   dSP_9_p;
  wire       [31:0]   dSP_10_p;
  wire       [31:0]   dSP_11_p;
  wire       [31:0]   dSP_12_p;
  wire       [31:0]   dSP_13_p;
  wire       [31:0]   dSP_14_p;
  wire       [31:0]   dSP_15_p;
  wire       [31:0]   dSP_16_p;
  wire       [31:0]   dSP_17_p;
  wire       [31:0]   dSP_18_p;
  wire       [31:0]   dSP_19_p;
  wire       [31:0]   dSP_20_p;
  wire       [31:0]   dSP_21_p;
  wire       [31:0]   dSP_22_p;
  wire       [31:0]   dSP_23_p;
  wire       [31:0]   dSP_24_p;
  wire       [31:0]   dSP_25_p;
  wire       [31:0]   dSP_26_p;
  wire       [31:0]   dSP_27_p;
  wire       [31:0]   dSP_28_p;
  wire       [31:0]   dSP_29_p;
  wire       [31:0]   dSP_30_p;
  wire       [31:0]   dSP_31_p;
  wire       [31:0]   dSP_32_p;
  wire       [31:0]   dSP_33_p;
  wire       [31:0]   dSP_34_p;
  wire       [31:0]   dSP_35_p;
  wire       [31:0]   dSP_36_p;
  wire       [31:0]   dSP_37_p;
  wire       [31:0]   dSP_38_p;
  wire       [31:0]   dSP_39_p;
  wire       [31:0]   dSP_40_p;
  wire       [31:0]   dSP_41_p;
  wire       [31:0]   dSP_42_p;
  wire       [31:0]   dSP_43_p;
  wire       [31:0]   dSP_44_p;
  wire       [31:0]   dSP_45_p;
  wire       [31:0]   dSP_46_p;
  wire       [31:0]   dSP_47_p;
  wire       [31:0]   dSP_48_p;
  wire       [31:0]   dSP_49_p;
  wire       [31:0]   dSP_50_p;
  wire       [31:0]   dSP_51_p;
  wire       [31:0]   dSP_52_p;
  wire       [31:0]   dSP_53_p;
  wire       [31:0]   dSP_54_p;
  wire       [31:0]   dSP_55_p;
  wire       [31:0]   dSP_56_p;
  wire       [31:0]   dSP_57_p;
  wire       [31:0]   dSP_58_p;
  wire       [31:0]   dSP_59_p;
  wire       [31:0]   dSP_60_p;
  wire       [31:0]   dSP_61_p;
  wire       [31:0]   dSP_62_p;
  wire       [31:0]   dSP_63_p;
  wire       [31:0]   dSP_64_p;
  wire       [31:0]   dSP_65_p;
  wire       [31:0]   dSP_66_p;
  wire       [31:0]   dSP_67_p;
  wire       [31:0]   dSP_68_p;
  wire       [31:0]   dSP_69_p;
  wire       [31:0]   dSP_70_p;
  wire       [31:0]   dSP_71_p;
  wire       [31:0]   dSP_72_p;
  wire       [31:0]   dSP_73_p;
  wire       [31:0]   dSP_74_p;
  wire       [31:0]   dSP_75_p;
  wire       [31:0]   dSP_76_p;
  wire       [31:0]   dSP_77_p;
  wire       [31:0]   dSP_78_p;
  wire       [31:0]   dSP_79_p;
  wire       [31:0]   dSP_80_p;
  wire       [31:0]   dSP_81_p;
  wire       [31:0]   dSP_82_p;
  wire       [31:0]   dSP_83_p;
  wire       [31:0]   dSP_84_p;
  wire       [31:0]   dSP_85_p;
  wire       [31:0]   dSP_86_p;
  wire       [31:0]   dSP_87_p;
  wire       [31:0]   dSP_88_p;
  wire       [31:0]   dSP_89_p;
  wire       [31:0]   dSP_90_p;
  wire       [31:0]   dSP_91_p;
  wire       [31:0]   dSP_92_p;
  wire       [31:0]   dSP_93_p;
  wire       [31:0]   dSP_94_p;
  wire       [31:0]   dSP_95_p;
  wire       [31:0]   dSP_96_p;
  wire       [31:0]   dSP_97_p;
  wire       [31:0]   dSP_98_p;
  wire       [31:0]   dSP_99_p;
  wire       [31:0]   dSP_100_p;
  wire       [31:0]   dSP_101_p;
  wire       [31:0]   dSP_102_p;
  wire       [31:0]   dSP_103_p;
  wire       [31:0]   dSP_104_p;
  wire       [31:0]   dSP_105_p;
  wire       [31:0]   dSP_106_p;
  wire       [31:0]   dSP_107_p;
  wire       [31:0]   dSP_108_p;
  wire       [31:0]   dSP_109_p;
  wire       [31:0]   dSP_110_p;
  wire       [31:0]   dSP_111_p;
  wire       [31:0]   dSP_112_p;
  wire       [31:0]   dSP_113_p;
  wire       [31:0]   dSP_114_p;
  wire       [31:0]   dSP_115_p;
  wire       [31:0]   dSP_116_p;
  wire       [31:0]   dSP_117_p;
  wire       [31:0]   dSP_118_p;
  wire       [31:0]   dSP_119_p;
  wire       [31:0]   dSP_120_p;
  wire       [31:0]   dSP_121_p;
  wire       [31:0]   dSP_122_p;
  wire       [31:0]   dSP_123_p;
  wire       [31:0]   dSP_124_p;
  wire       [31:0]   dSP_125_p;
  wire       [31:0]   dSP_126_p;
  wire       [31:0]   dSP_127_p;
  wire       [31:0]   dSP_128_p;
  wire       [31:0]   dSP_129_p;
  wire       [31:0]   dSP_130_p;
  wire       [31:0]   dSP_131_p;
  wire       [31:0]   dSP_132_p;
  wire       [31:0]   dSP_133_p;
  wire       [31:0]   dSP_134_p;
  wire       [31:0]   dSP_135_p;
  wire       [31:0]   dSP_136_p;
  wire       [31:0]   dSP_137_p;
  wire       [31:0]   dSP_138_p;
  wire       [31:0]   dSP_139_p;
  wire       [31:0]   dSP_140_p;
  wire       [31:0]   dSP_141_p;
  wire       [31:0]   dSP_142_p;
  wire       [31:0]   dSP_143_p;
  wire       [31:0]   dSP_144_p;
  wire       [31:0]   dSP_145_p;
  wire       [31:0]   dSP_146_p;
  wire       [31:0]   dSP_147_p;
  wire       [31:0]   dSP_148_p;
  wire       [31:0]   dSP_149_p;
  wire       [31:0]   dSP_150_p;
  wire       [31:0]   dSP_151_p;
  wire       [31:0]   dSP_152_p;
  wire       [31:0]   dSP_153_p;
  wire       [31:0]   dSP_154_p;
  wire       [31:0]   dSP_155_p;
  wire       [31:0]   dSP_156_p;
  wire       [31:0]   dSP_157_p;
  wire       [31:0]   dSP_158_p;
  wire       [31:0]   dSP_159_p;
  wire       [31:0]   dSP_160_p;
  wire       [31:0]   dSP_161_p;
  wire       [31:0]   dSP_162_p;
  wire       [31:0]   dSP_163_p;
  wire       [31:0]   dSP_164_p;
  wire       [31:0]   dSP_165_p;
  wire       [31:0]   dSP_166_p;
  wire       [31:0]   dSP_167_p;
  wire       [31:0]   dSP_168_p;
  wire       [31:0]   dSP_169_p;
  wire       [31:0]   dSP_170_p;
  wire       [31:0]   dSP_171_p;
  wire       [31:0]   dSP_172_p;
  wire       [31:0]   dSP_173_p;
  wire       [31:0]   dSP_174_p;
  wire       [31:0]   dSP_175_p;
  wire       [31:0]   dSP_176_p;
  wire       [31:0]   dSP_177_p;
  wire       [31:0]   dSP_178_p;
  wire       [31:0]   dSP_179_p;
  wire       [31:0]   dSP_180_p;
  wire       [31:0]   dSP_181_p;
  wire       [31:0]   dSP_182_p;
  wire       [31:0]   dSP_183_p;
  wire       [31:0]   dSP_184_p;
  wire       [31:0]   dSP_185_p;
  wire       [31:0]   dSP_186_p;
  wire       [31:0]   dSP_187_p;
  wire       [31:0]   dSP_188_p;
  wire       [31:0]   dSP_189_p;
  wire       [31:0]   dSP_190_p;
  wire       [31:0]   dSP_191_p;
  wire       [31:0]   dSP_192_p;
  wire       [31:0]   dSP_193_p;
  wire       [31:0]   dSP_194_p;
  wire       [31:0]   dSP_195_p;
  wire       [31:0]   dSP_196_p;
  wire       [31:0]   dSP_197_p;
  wire       [31:0]   dSP_198_p;
  wire       [31:0]   dSP_199_p;
  wire       [31:0]   dSP_200_p;
  wire       [31:0]   dSP_201_p;
  wire       [31:0]   dSP_202_p;
  wire       [31:0]   dSP_203_p;
  wire       [31:0]   dSP_204_p;
  wire       [31:0]   dSP_205_p;
  wire       [31:0]   dSP_206_p;
  wire       [31:0]   dSP_207_p;
  wire       [31:0]   dSP_208_p;
  wire       [31:0]   dSP_209_p;
  wire       [31:0]   dSP_210_p;
  wire       [31:0]   dSP_211_p;
  wire       [31:0]   dSP_212_p;
  wire       [31:0]   dSP_213_p;
  wire       [31:0]   dSP_214_p;
  wire       [31:0]   dSP_215_p;
  wire       [31:0]   dSP_216_p;
  wire       [31:0]   dSP_217_p;
  wire       [31:0]   dSP_218_p;
  wire       [31:0]   dSP_219_p;
  wire       [31:0]   dSP_220_p;
  wire       [31:0]   dSP_221_p;
  wire       [31:0]   dSP_222_p;
  wire       [31:0]   dSP_223_p;
  wire       [31:0]   dSP_224_p;
  wire       [31:0]   dSP_225_p;
  wire       [31:0]   dSP_226_p;
  wire       [31:0]   dSP_227_p;
  wire       [31:0]   dSP_228_p;
  wire       [31:0]   dSP_229_p;
  wire       [31:0]   dSP_230_p;
  wire       [31:0]   dSP_231_p;
  wire       [31:0]   dSP_232_p;
  wire       [31:0]   dSP_233_p;
  wire       [31:0]   dSP_234_p;
  wire       [31:0]   dSP_235_p;
  wire       [31:0]   dSP_236_p;
  wire       [31:0]   dSP_237_p;
  wire       [31:0]   dSP_238_p;
  wire       [31:0]   dSP_239_p;
  wire       [31:0]   dSP_240_p;
  wire       [31:0]   dSP_241_p;
  wire       [31:0]   dSP_242_p;
  wire       [31:0]   dSP_243_p;
  wire       [31:0]   dSP_244_p;
  wire       [31:0]   dSP_245_p;
  wire       [31:0]   dSP_246_p;
  wire       [31:0]   dSP_247_p;
  wire       [31:0]   dSP_248_p;
  wire       [31:0]   dSP_249_p;
  wire       [31:0]   dSP_250_p;
  wire       [31:0]   dSP_251_p;
  wire       [31:0]   dSP_252_p;
  wire       [31:0]   dSP_253_p;
  wire       [31:0]   dSP_254_p;
  wire       [31:0]   dSP_255_p;
  wire       [31:0]   dSP_256_p;
  wire       [31:0]   dSP_257_p;
  wire       [31:0]   dSP_258_p;
  wire       [31:0]   dSP_259_p;
  wire       [31:0]   dSP_260_p;
  wire       [31:0]   dSP_261_p;
  wire       [31:0]   dSP_262_p;
  wire       [31:0]   dSP_263_p;
  wire       [31:0]   dSP_264_p;
  wire       [31:0]   dSP_265_p;
  wire       [31:0]   dSP_266_p;
  wire       [31:0]   dSP_267_p;
  wire       [31:0]   dSP_268_p;
  wire       [31:0]   dSP_269_p;
  wire       [31:0]   dSP_270_p;
  wire       [31:0]   dSP_271_p;
  wire       [31:0]   dSP_272_p;
  wire       [31:0]   dSP_273_p;
  wire       [31:0]   dSP_274_p;
  wire       [31:0]   dSP_275_p;
  wire       [31:0]   dSP_276_p;
  wire       [31:0]   dSP_277_p;
  wire       [31:0]   dSP_278_p;
  wire       [31:0]   dSP_279_p;
  wire       [31:0]   dSP_280_p;
  wire       [31:0]   dSP_281_p;
  wire       [31:0]   dSP_282_p;
  wire       [31:0]   dSP_283_p;
  wire       [31:0]   dSP_284_p;
  wire       [31:0]   dSP_285_p;
  wire       [31:0]   dSP_286_p;
  wire       [31:0]   dSP_287_p;
  wire       [31:0]   dSP_288_p;
  wire       [31:0]   dSP_289_p;
  wire       [31:0]   dSP_290_p;
  wire       [31:0]   dSP_291_p;
  wire       [31:0]   dSP_292_p;
  wire       [31:0]   dSP_293_p;
  wire       [31:0]   dSP_294_p;
  wire       [31:0]   dSP_295_p;
  wire       [31:0]   dSP_296_p;
  wire       [31:0]   dSP_297_p;
  wire       [31:0]   dSP_298_p;
  wire       [31:0]   dSP_299_p;
  wire       [31:0]   dSP_300_p;
  wire       [31:0]   dSP_301_p;
  wire       [31:0]   dSP_302_p;
  wire       [31:0]   dSP_303_p;
  wire       [31:0]   dSP_304_p;
  wire       [31:0]   dSP_305_p;
  wire       [31:0]   dSP_306_p;
  wire       [31:0]   dSP_307_p;
  wire       [31:0]   dSP_308_p;
  wire       [31:0]   dSP_309_p;
  wire       [31:0]   dSP_310_p;
  wire       [31:0]   dSP_311_p;
  wire       [31:0]   dSP_312_p;
  wire       [31:0]   dSP_313_p;
  wire       [31:0]   dSP_314_p;
  wire       [31:0]   dSP_315_p;
  wire       [31:0]   dSP_316_p;
  wire       [31:0]   dSP_317_p;
  wire       [31:0]   dSP_318_p;
  wire       [31:0]   dSP_319_p;
  wire       [31:0]   dSP_320_p;
  wire       [31:0]   dSP_321_p;
  wire       [31:0]   dSP_322_p;
  wire       [31:0]   dSP_323_p;
  wire       [31:0]   dSP_324_p;
  wire       [31:0]   dSP_325_p;
  wire       [31:0]   dSP_326_p;
  wire       [31:0]   dSP_327_p;
  wire       [31:0]   dSP_328_p;
  wire       [31:0]   dSP_329_p;
  wire       [31:0]   dSP_330_p;
  wire       [31:0]   dSP_331_p;
  wire       [31:0]   dSP_332_p;
  wire       [31:0]   dSP_333_p;
  wire       [31:0]   dSP_334_p;
  wire       [31:0]   dSP_335_p;
  wire       [31:0]   dSP_336_p;
  wire       [31:0]   dSP_337_p;
  wire       [31:0]   dSP_338_p;
  wire       [31:0]   dSP_339_p;
  wire       [31:0]   dSP_340_p;
  wire       [31:0]   dSP_341_p;
  wire       [31:0]   dSP_342_p;
  wire       [31:0]   dSP_343_p;
  wire       [31:0]   dSP_344_p;
  wire       [31:0]   dSP_345_p;
  wire       [31:0]   dSP_346_p;
  wire       [31:0]   dSP_347_p;
  wire       [31:0]   dSP_348_p;
  wire       [31:0]   dSP_349_p;
  wire       [31:0]   dSP_350_p;
  wire       [31:0]   dSP_351_p;
  wire       [31:0]   dSP_352_p;
  wire       [31:0]   dSP_353_p;
  wire       [31:0]   dSP_354_p;
  wire       [31:0]   dSP_355_p;
  wire       [31:0]   dSP_356_p;
  wire       [31:0]   dSP_357_p;
  wire       [31:0]   dSP_358_p;
  wire       [31:0]   dSP_359_p;
  wire       [31:0]   dSP_360_p;
  wire       [31:0]   dSP_361_p;
  wire       [31:0]   dSP_362_p;
  wire       [31:0]   dSP_363_p;
  wire       [31:0]   dSP_364_p;
  wire       [31:0]   dSP_365_p;
  wire       [31:0]   dSP_366_p;
  wire       [31:0]   dSP_367_p;
  wire       [31:0]   dSP_368_p;
  wire       [31:0]   dSP_369_p;
  wire       [31:0]   dSP_370_p;
  wire       [31:0]   dSP_371_p;
  wire       [31:0]   dSP_372_p;
  wire       [31:0]   dSP_373_p;
  wire       [31:0]   dSP_374_p;
  wire       [31:0]   dSP_375_p;
  wire       [31:0]   dSP_376_p;
  wire       [31:0]   dSP_377_p;
  wire       [31:0]   dSP_378_p;
  wire       [31:0]   dSP_379_p;
  wire       [31:0]   dSP_380_p;
  wire       [31:0]   dSP_381_p;
  wire       [31:0]   dSP_382_p;
  wire       [31:0]   dSP_383_p;
  wire       [31:0]   dSP_384_p;
  wire       [31:0]   dSP_385_p;
  wire       [31:0]   dSP_386_p;
  wire       [31:0]   dSP_387_p;
  wire       [31:0]   dSP_388_p;
  wire       [31:0]   dSP_389_p;
  wire       [31:0]   dSP_390_p;
  wire       [31:0]   dSP_391_p;
  wire       [31:0]   dSP_392_p;
  wire       [31:0]   dSP_393_p;
  wire       [31:0]   dSP_394_p;
  wire       [31:0]   dSP_395_p;
  wire       [31:0]   dSP_396_p;
  wire       [31:0]   dSP_397_p;
  wire       [31:0]   dSP_398_p;
  wire       [31:0]   dSP_399_p;
  wire       [31:0]   dSP_400_p;
  wire       [31:0]   dSP_401_p;
  wire       [31:0]   dSP_402_p;
  wire       [31:0]   dSP_403_p;
  wire       [31:0]   dSP_404_p;
  wire       [31:0]   dSP_405_p;
  wire       [31:0]   dSP_406_p;
  wire       [31:0]   dSP_407_p;
  wire       [31:0]   dSP_408_p;
  wire       [31:0]   dSP_409_p;
  wire       [31:0]   dSP_410_p;
  wire       [31:0]   dSP_411_p;
  wire       [31:0]   dSP_412_p;
  wire       [31:0]   dSP_413_p;
  wire       [31:0]   dSP_414_p;
  wire       [31:0]   dSP_415_p;
  wire       [31:0]   dSP_416_p;
  wire       [31:0]   dSP_417_p;
  wire       [31:0]   dSP_418_p;
  wire       [31:0]   dSP_419_p;
  wire       [31:0]   dSP_420_p;
  wire       [31:0]   dSP_421_p;
  wire       [31:0]   dSP_422_p;
  wire       [31:0]   dSP_423_p;
  wire       [31:0]   dSP_424_p;
  wire       [31:0]   dSP_425_p;
  wire       [31:0]   dSP_426_p;
  wire       [31:0]   dSP_427_p;
  wire       [31:0]   dSP_428_p;
  wire       [31:0]   dSP_429_p;
  wire       [31:0]   dSP_430_p;
  wire       [31:0]   dSP_431_p;
  wire       [31:0]   dSP_432_p;
  wire       [31:0]   dSP_433_p;
  wire       [31:0]   dSP_434_p;
  wire       [31:0]   dSP_435_p;
  wire       [31:0]   dSP_436_p;
  wire       [31:0]   dSP_437_p;
  wire       [31:0]   dSP_438_p;
  wire       [31:0]   dSP_439_p;
  wire       [31:0]   dSP_440_p;
  wire       [31:0]   dSP_441_p;
  wire       [31:0]   dSP_442_p;
  wire       [31:0]   dSP_443_p;
  wire       [31:0]   dSP_444_p;
  wire       [31:0]   dSP_445_p;
  wire       [31:0]   dSP_446_p;
  wire       [31:0]   dSP_447_p;
  wire       [31:0]   dSP_448_p;
  wire       [31:0]   dSP_449_p;
  wire       [31:0]   dSP_450_p;
  wire       [31:0]   dSP_451_p;
  wire       [31:0]   dSP_452_p;
  wire       [31:0]   dSP_453_p;
  wire       [31:0]   dSP_454_p;
  wire       [31:0]   dSP_455_p;
  wire       [31:0]   dSP_456_p;
  wire       [31:0]   dSP_457_p;
  wire       [31:0]   dSP_458_p;
  wire       [31:0]   dSP_459_p;
  wire       [31:0]   dSP_460_p;
  wire       [31:0]   dSP_461_p;
  wire       [31:0]   dSP_462_p;
  wire       [31:0]   dSP_463_p;
  wire       [31:0]   dSP_464_p;
  wire       [31:0]   dSP_465_p;
  wire       [31:0]   dSP_466_p;
  wire       [31:0]   dSP_467_p;
  wire       [31:0]   dSP_468_p;
  wire       [31:0]   dSP_469_p;
  wire       [31:0]   dSP_470_p;
  wire       [31:0]   dSP_471_p;
  wire       [31:0]   dSP_472_p;
  wire       [31:0]   dSP_473_p;
  wire       [31:0]   dSP_474_p;
  wire       [31:0]   dSP_475_p;
  wire       [31:0]   dSP_476_p;
  wire       [31:0]   dSP_477_p;
  wire       [31:0]   dSP_478_p;
  wire       [31:0]   dSP_479_p;
  wire       [31:0]   dSP_480_p;
  wire       [31:0]   dSP_481_p;
  wire       [31:0]   dSP_482_p;
  wire       [31:0]   dSP_483_p;
  wire       [31:0]   dSP_484_p;
  wire       [31:0]   dSP_485_p;
  wire       [31:0]   dSP_486_p;
  wire       [31:0]   dSP_487_p;
  wire       [31:0]   dSP_488_p;
  wire       [31:0]   dSP_489_p;
  wire       [31:0]   dSP_490_p;
  wire       [31:0]   dSP_491_p;
  wire       [31:0]   dSP_492_p;
  wire       [31:0]   dSP_493_p;
  wire       [31:0]   dSP_494_p;
  wire       [31:0]   dSP_495_p;
  wire       [31:0]   dSP_496_p;
  wire       [31:0]   dSP_497_p;
  wire       [31:0]   dSP_498_p;
  wire       [31:0]   dSP_499_p;
  wire       [31:0]   dSP_500_p;
  wire       [31:0]   dSP_501_p;
  wire       [31:0]   dSP_502_p;
  wire       [31:0]   dSP_503_p;
  wire       [31:0]   dSP_504_p;
  wire       [31:0]   dSP_505_p;
  wire       [31:0]   dSP_506_p;
  wire       [31:0]   dSP_507_p;
  wire       [31:0]   dSP_508_p;
  wire       [31:0]   dSP_509_p;
  wire       [31:0]   dSP_510_p;
  wire       [31:0]   dSP_511_p;
  wire       [31:0]   dSP_512_p;
  wire       [31:0]   dSP_513_p;
  wire       [31:0]   dSP_514_p;
  wire       [31:0]   dSP_515_p;
  wire       [31:0]   dSP_516_p;
  wire       [31:0]   dSP_517_p;
  wire       [31:0]   dSP_518_p;
  wire       [31:0]   dSP_519_p;
  wire       [31:0]   dSP_520_p;
  wire       [31:0]   dSP_521_p;
  wire       [31:0]   dSP_522_p;
  wire       [31:0]   dSP_523_p;
  wire       [31:0]   dSP_524_p;
  wire       [31:0]   dSP_525_p;
  wire       [31:0]   dSP_526_p;
  wire       [31:0]   dSP_527_p;
  wire       [31:0]   dSP_528_p;
  wire       [31:0]   dSP_529_p;
  wire       [31:0]   dSP_530_p;
  wire       [31:0]   dSP_531_p;
  wire       [31:0]   dSP_532_p;
  wire       [31:0]   dSP_533_p;
  wire       [31:0]   dSP_534_p;
  wire       [31:0]   dSP_535_p;
  wire       [31:0]   dSP_536_p;
  wire       [31:0]   dSP_537_p;
  wire       [31:0]   dSP_538_p;
  wire       [31:0]   dSP_539_p;
  wire       [31:0]   dSP_540_p;
  wire       [31:0]   dSP_541_p;
  wire       [31:0]   dSP_542_p;
  wire       [31:0]   dSP_543_p;
  wire       [31:0]   dSP_544_p;
  wire       [31:0]   dSP_545_p;
  wire       [31:0]   dSP_546_p;
  wire       [31:0]   dSP_547_p;
  wire       [31:0]   dSP_548_p;
  wire       [31:0]   dSP_549_p;
  wire       [31:0]   dSP_550_p;
  wire       [31:0]   dSP_551_p;
  wire       [31:0]   dSP_552_p;
  wire       [31:0]   dSP_553_p;
  wire       [31:0]   dSP_554_p;
  wire       [31:0]   dSP_555_p;
  wire       [31:0]   dSP_556_p;
  wire       [31:0]   dSP_557_p;
  wire       [31:0]   dSP_558_p;
  wire       [31:0]   dSP_559_p;
  wire       [31:0]   dSP_560_p;
  wire       [31:0]   dSP_561_p;
  wire       [31:0]   dSP_562_p;
  wire       [31:0]   dSP_563_p;
  wire       [31:0]   dSP_564_p;
  wire       [31:0]   dSP_565_p;
  wire       [31:0]   dSP_566_p;
  wire       [31:0]   dSP_567_p;
  wire       [31:0]   dSP_568_p;
  wire       [31:0]   dSP_569_p;
  wire       [31:0]   dSP_570_p;
  wire       [31:0]   dSP_571_p;
  wire       [31:0]   dSP_572_p;
  wire       [31:0]   dSP_573_p;
  wire       [31:0]   dSP_574_p;
  wire       [31:0]   dSP_575_p;
  wire       [31:0]   dSP_576_p;
  wire       [31:0]   dSP_577_p;
  wire       [31:0]   dSP_578_p;
  wire       [31:0]   dSP_579_p;
  wire       [31:0]   dSP_580_p;
  wire       [31:0]   dSP_581_p;
  wire       [31:0]   dSP_582_p;
  wire       [31:0]   dSP_583_p;
  wire       [31:0]   dSP_584_p;
  wire       [31:0]   dSP_585_p;
  wire       [31:0]   dSP_586_p;
  wire       [31:0]   dSP_587_p;
  wire       [31:0]   dSP_588_p;
  wire       [31:0]   dSP_589_p;
  wire       [31:0]   dSP_590_p;
  wire       [31:0]   dSP_591_p;
  wire       [31:0]   dSP_592_p;
  wire       [31:0]   dSP_593_p;
  wire       [31:0]   dSP_594_p;
  wire       [31:0]   dSP_595_p;
  wire       [31:0]   dSP_596_p;
  wire       [31:0]   dSP_597_p;
  wire       [31:0]   dSP_598_p;
  wire       [31:0]   dSP_599_p;
  wire       [31:0]   dSP_600_p;
  wire       [31:0]   dSP_601_p;
  wire       [31:0]   dSP_602_p;
  wire       [31:0]   dSP_603_p;
  wire       [31:0]   dSP_604_p;
  wire       [31:0]   dSP_605_p;
  wire       [31:0]   dSP_606_p;
  wire       [31:0]   dSP_607_p;
  wire       [31:0]   dSP_608_p;
  wire       [31:0]   dSP_609_p;
  wire       [31:0]   dSP_610_p;
  wire       [31:0]   dSP_611_p;
  wire       [31:0]   dSP_612_p;
  wire       [31:0]   dSP_613_p;
  wire       [31:0]   dSP_614_p;
  wire       [31:0]   dSP_615_p;
  wire       [31:0]   dSP_616_p;
  wire       [31:0]   dSP_617_p;
  wire       [31:0]   dSP_618_p;
  wire       [31:0]   dSP_619_p;
  wire       [31:0]   dSP_620_p;
  wire       [31:0]   dSP_621_p;
  wire       [31:0]   dSP_622_p;
  wire       [31:0]   dSP_623_p;
  wire       [31:0]   dSP_624_p;
  wire       [31:0]   dSP_625_p;
  wire       [31:0]   dSP_626_p;
  wire       [31:0]   dSP_627_p;
  wire       [31:0]   dSP_628_p;
  wire       [31:0]   dSP_629_p;
  wire       [31:0]   dSP_630_p;
  wire       [31:0]   dSP_631_p;
  wire       [31:0]   dSP_632_p;
  wire       [31:0]   dSP_633_p;
  wire       [31:0]   dSP_634_p;
  wire       [31:0]   dSP_635_p;
  wire       [31:0]   dSP_636_p;
  wire       [31:0]   dSP_637_p;
  wire       [31:0]   dSP_638_p;
  wire       [31:0]   dSP_639_p;
  wire       [31:0]   dSP_640_p;
  wire       [31:0]   dSP_641_p;
  wire       [31:0]   dSP_642_p;
  wire       [31:0]   dSP_643_p;
  wire       [31:0]   dSP_644_p;
  wire       [31:0]   dSP_645_p;
  wire       [31:0]   dSP_646_p;
  wire       [31:0]   dSP_647_p;
  wire       [31:0]   dSP_648_p;
  wire       [31:0]   dSP_649_p;
  wire       [31:0]   dSP_650_p;
  wire       [31:0]   dSP_651_p;
  wire       [31:0]   dSP_652_p;
  wire       [31:0]   dSP_653_p;
  wire       [31:0]   dSP_654_p;
  wire       [31:0]   dSP_655_p;
  wire       [31:0]   dSP_656_p;
  wire       [31:0]   dSP_657_p;
  wire       [31:0]   dSP_658_p;
  wire       [31:0]   dSP_659_p;
  wire       [31:0]   dSP_660_p;
  wire       [31:0]   dSP_661_p;
  wire       [31:0]   dSP_662_p;
  wire       [31:0]   dSP_663_p;
  wire       [31:0]   dSP_664_p;
  wire       [31:0]   dSP_665_p;
  wire       [31:0]   dSP_666_p;
  wire       [31:0]   dSP_667_p;
  wire       [31:0]   dSP_668_p;
  wire       [31:0]   dSP_669_p;
  wire       [31:0]   dSP_670_p;
  wire       [31:0]   dSP_671_p;
  wire       [31:0]   dSP_672_p;
  wire       [31:0]   dSP_673_p;
  wire       [31:0]   dSP_674_p;
  wire       [31:0]   dSP_675_p;
  wire       [31:0]   dSP_676_p;
  wire       [31:0]   dSP_677_p;
  wire       [31:0]   dSP_678_p;
  wire       [31:0]   dSP_679_p;
  wire       [31:0]   dSP_680_p;
  wire       [31:0]   dSP_681_p;
  wire       [31:0]   dSP_682_p;
  wire       [31:0]   dSP_683_p;
  wire       [31:0]   dSP_684_p;
  wire       [31:0]   dSP_685_p;
  wire       [31:0]   dSP_686_p;
  wire       [31:0]   dSP_687_p;
  wire       [31:0]   dSP_688_p;
  wire       [31:0]   dSP_689_p;
  wire       [31:0]   dSP_690_p;
  wire       [31:0]   dSP_691_p;
  wire       [31:0]   dSP_692_p;
  wire       [31:0]   dSP_693_p;
  wire       [31:0]   dSP_694_p;
  wire       [31:0]   dSP_695_p;
  wire       [31:0]   dSP_696_p;
  wire       [31:0]   dSP_697_p;
  wire       [31:0]   dSP_698_p;
  wire       [31:0]   dSP_699_p;
  wire       [31:0]   dSP_700_p;
  wire       [31:0]   dSP_701_p;
  wire       [31:0]   dSP_702_p;
  wire       [31:0]   dSP_703_p;
  wire       [31:0]   dSP_704_p;
  wire       [31:0]   dSP_705_p;
  wire       [31:0]   dSP_706_p;
  wire       [31:0]   dSP_707_p;
  wire       [31:0]   dSP_708_p;
  wire       [31:0]   dSP_709_p;
  wire       [31:0]   dSP_710_p;
  wire       [31:0]   dSP_711_p;
  wire       [31:0]   dSP_712_p;
  wire       [31:0]   dSP_713_p;
  wire       [31:0]   dSP_714_p;
  wire       [31:0]   dSP_715_p;
  wire       [31:0]   dSP_716_p;
  wire       [31:0]   dSP_717_p;
  wire       [31:0]   dSP_718_p;
  wire       [31:0]   dSP_719_p;
  wire       [31:0]   dSP_720_p;
  wire       [31:0]   dSP_721_p;
  wire       [31:0]   dSP_722_p;
  wire       [31:0]   dSP_723_p;
  wire       [31:0]   dSP_724_p;
  wire       [31:0]   dSP_725_p;
  wire       [31:0]   dSP_726_p;
  wire       [31:0]   dSP_727_p;
  wire       [31:0]   dSP_728_p;
  wire       [31:0]   dSP_729_p;
  wire       [31:0]   dSP_730_p;
  wire       [31:0]   dSP_731_p;
  wire       [31:0]   dSP_732_p;
  wire       [31:0]   dSP_733_p;
  wire       [31:0]   dSP_734_p;
  wire       [31:0]   dSP_735_p;
  wire       [31:0]   dSP_736_p;
  wire       [31:0]   dSP_737_p;
  wire       [31:0]   dSP_738_p;
  wire       [31:0]   dSP_739_p;
  wire       [31:0]   dSP_740_p;
  wire       [31:0]   dSP_741_p;
  wire       [31:0]   dSP_742_p;
  wire       [31:0]   dSP_743_p;
  wire       [31:0]   dSP_744_p;
  wire       [31:0]   dSP_745_p;
  wire       [31:0]   dSP_746_p;
  wire       [31:0]   dSP_747_p;
  wire       [31:0]   dSP_748_p;
  wire       [31:0]   dSP_749_p;
  wire       [31:0]   dSP_750_p;
  wire       [31:0]   dSP_751_p;
  wire       [31:0]   dSP_752_p;
  wire       [31:0]   dSP_753_p;
  wire       [31:0]   dSP_754_p;
  wire       [31:0]   dSP_755_p;
  wire       [31:0]   dSP_756_p;
  wire       [31:0]   dSP_757_p;
  wire       [31:0]   dSP_758_p;
  wire       [31:0]   dSP_759_p;
  wire       [31:0]   dSP_760_p;
  wire       [31:0]   dSP_761_p;
  wire       [31:0]   dSP_762_p;
  wire       [31:0]   dSP_763_p;
  wire       [31:0]   dSP_764_p;
  wire       [31:0]   dSP_765_p;
  wire       [31:0]   dSP_766_p;
  wire       [31:0]   dSP_767_p;
  wire       [31:0]   dSP_768_p;
  wire       [31:0]   dSP_769_p;
  wire       [31:0]   dSP_770_p;
  wire       [31:0]   dSP_771_p;
  wire       [31:0]   dSP_772_p;
  wire       [31:0]   dSP_773_p;
  wire       [31:0]   dSP_774_p;
  wire       [31:0]   dSP_775_p;
  wire       [31:0]   dSP_776_p;
  wire       [31:0]   dSP_777_p;
  wire       [31:0]   dSP_778_p;
  wire       [31:0]   dSP_779_p;
  wire       [31:0]   dSP_780_p;
  wire       [31:0]   dSP_781_p;
  wire       [31:0]   dSP_782_p;
  wire       [31:0]   dSP_783_p;
  wire       [31:0]   dSP_784_p;
  wire       [31:0]   dSP_785_p;
  wire       [31:0]   dSP_786_p;
  wire       [31:0]   dSP_787_p;
  wire       [31:0]   dSP_788_p;
  wire       [31:0]   dSP_789_p;
  wire       [31:0]   dSP_790_p;
  wire       [31:0]   dSP_791_p;
  wire       [31:0]   dSP_792_p;
  wire       [31:0]   dSP_793_p;
  wire       [31:0]   dSP_794_p;
  wire       [31:0]   dSP_795_p;
  wire       [31:0]   dSP_796_p;
  wire       [31:0]   dSP_797_p;
  wire       [31:0]   dSP_798_p;
  wire       [31:0]   dSP_799_p;
  wire       [31:0]   dSP_800_p;
  wire       [31:0]   dSP_801_p;
  wire       [31:0]   dSP_802_p;
  wire       [31:0]   dSP_803_p;
  wire       [31:0]   dSP_804_p;
  wire       [31:0]   dSP_805_p;
  wire       [31:0]   dSP_806_p;
  wire       [31:0]   dSP_807_p;
  wire       [31:0]   dSP_808_p;
  wire       [31:0]   dSP_809_p;
  wire       [31:0]   dSP_810_p;
  wire       [31:0]   dSP_811_p;
  wire       [31:0]   dSP_812_p;
  wire       [31:0]   dSP_813_p;
  wire       [31:0]   dSP_814_p;
  wire       [31:0]   dSP_815_p;
  wire       [31:0]   dSP_816_p;
  wire       [31:0]   dSP_817_p;
  wire       [31:0]   dSP_818_p;
  wire       [31:0]   dSP_819_p;
  wire       [31:0]   dSP_820_p;
  wire       [31:0]   dSP_821_p;
  wire       [31:0]   dSP_822_p;
  wire       [31:0]   dSP_823_p;
  wire       [31:0]   dSP_824_p;
  wire       [31:0]   dSP_825_p;
  wire       [31:0]   dSP_826_p;
  wire       [31:0]   dSP_827_p;
  wire       [31:0]   dSP_828_p;
  wire       [31:0]   dSP_829_p;
  wire       [31:0]   dSP_830_p;
  wire       [31:0]   dSP_831_p;
  wire       [31:0]   dSP_832_p;
  wire       [31:0]   dSP_833_p;
  wire       [31:0]   dSP_834_p;
  wire       [31:0]   dSP_835_p;
  wire       [31:0]   dSP_836_p;
  wire       [31:0]   dSP_837_p;
  wire       [31:0]   dSP_838_p;
  wire       [31:0]   dSP_839_p;
  wire       [31:0]   dSP_840_p;
  wire       [31:0]   dSP_841_p;
  wire       [31:0]   dSP_842_p;
  wire       [31:0]   dSP_843_p;
  wire       [31:0]   dSP_844_p;
  wire       [31:0]   dSP_845_p;
  wire       [31:0]   dSP_846_p;
  wire       [31:0]   dSP_847_p;
  wire       [31:0]   dSP_848_p;
  wire       [31:0]   dSP_849_p;
  wire       [31:0]   dSP_850_p;
  wire       [31:0]   dSP_851_p;
  wire       [31:0]   dSP_852_p;
  wire       [31:0]   dSP_853_p;
  wire       [31:0]   dSP_854_p;
  wire       [31:0]   dSP_855_p;
  wire       [31:0]   dSP_856_p;
  wire       [31:0]   dSP_857_p;
  wire       [31:0]   dSP_858_p;
  wire       [31:0]   dSP_859_p;
  wire       [31:0]   dSP_860_p;
  wire       [31:0]   dSP_861_p;
  wire       [31:0]   dSP_862_p;
  wire       [31:0]   dSP_863_p;
  wire       [31:0]   dSP_864_p;
  wire       [31:0]   dSP_865_p;
  wire       [31:0]   dSP_866_p;
  wire       [31:0]   dSP_867_p;
  wire       [31:0]   dSP_868_p;
  wire       [31:0]   dSP_869_p;
  wire       [31:0]   dSP_870_p;
  wire       [31:0]   dSP_871_p;
  wire       [31:0]   dSP_872_p;
  wire       [31:0]   dSP_873_p;
  wire       [31:0]   dSP_874_p;
  wire       [31:0]   dSP_875_p;
  wire       [31:0]   dSP_876_p;
  wire       [31:0]   dSP_877_p;
  wire       [31:0]   dSP_878_p;
  wire       [31:0]   dSP_879_p;
  wire       [31:0]   dSP_880_p;
  wire       [31:0]   dSP_881_p;
  wire       [31:0]   dSP_882_p;
  wire       [31:0]   dSP_883_p;
  wire       [31:0]   dSP_884_p;
  wire       [31:0]   dSP_885_p;
  wire       [31:0]   dSP_886_p;
  wire       [31:0]   dSP_887_p;
  wire       [31:0]   dSP_888_p;
  wire       [31:0]   dSP_889_p;
  wire       [31:0]   dSP_890_p;
  wire       [31:0]   dSP_891_p;
  wire       [31:0]   dSP_892_p;
  wire       [31:0]   dSP_893_p;
  wire       [31:0]   dSP_894_p;
  wire       [31:0]   dSP_895_p;
  wire       [31:0]   dSP_896_p;
  wire       [31:0]   dSP_897_p;
  wire       [31:0]   dSP_898_p;
  wire       [31:0]   dSP_899_p;
  wire       [31:0]   dSP_900_p;
  wire       [31:0]   dSP_901_p;
  wire       [31:0]   dSP_902_p;
  wire       [31:0]   dSP_903_p;
  wire       [31:0]   dSP_904_p;
  wire       [31:0]   dSP_905_p;
  wire       [31:0]   dSP_906_p;
  wire       [31:0]   dSP_907_p;
  wire       [31:0]   dSP_908_p;
  wire       [31:0]   dSP_909_p;
  wire       [31:0]   dSP_910_p;
  wire       [31:0]   dSP_911_p;
  wire       [31:0]   dSP_912_p;
  wire       [31:0]   dSP_913_p;
  wire       [31:0]   dSP_914_p;
  wire       [31:0]   dSP_915_p;
  wire       [31:0]   dSP_916_p;
  wire       [31:0]   dSP_917_p;
  wire       [31:0]   dSP_918_p;
  wire       [31:0]   dSP_919_p;
  wire       [31:0]   dSP_920_p;
  wire       [31:0]   dSP_921_p;
  wire       [31:0]   dSP_922_p;
  wire       [31:0]   dSP_923_p;
  wire       [31:0]   dSP_924_p;
  wire       [31:0]   dSP_925_p;
  wire       [31:0]   dSP_926_p;
  wire       [31:0]   dSP_927_p;
  wire       [31:0]   dSP_928_p;
  wire       [31:0]   dSP_929_p;
  wire       [31:0]   dSP_930_p;
  wire       [31:0]   dSP_931_p;
  wire       [31:0]   dSP_932_p;
  wire       [31:0]   dSP_933_p;
  wire       [31:0]   dSP_934_p;
  wire       [31:0]   dSP_935_p;
  wire       [31:0]   dSP_936_p;
  wire       [31:0]   dSP_937_p;
  wire       [31:0]   dSP_938_p;
  wire       [31:0]   dSP_939_p;
  wire       [31:0]   dSP_940_p;
  wire       [31:0]   dSP_941_p;
  wire       [31:0]   dSP_942_p;
  wire       [31:0]   dSP_943_p;
  wire       [31:0]   dSP_944_p;
  wire       [31:0]   dSP_945_p;
  wire       [31:0]   dSP_946_p;
  wire       [31:0]   dSP_947_p;
  wire       [31:0]   dSP_948_p;
  wire       [31:0]   dSP_949_p;
  wire       [31:0]   dSP_950_p;
  wire       [31:0]   dSP_951_p;
  wire       [31:0]   dSP_952_p;
  wire       [31:0]   dSP_953_p;
  wire       [31:0]   dSP_954_p;
  wire       [31:0]   dSP_955_p;
  wire       [31:0]   dSP_956_p;
  wire       [31:0]   dSP_957_p;
  wire       [31:0]   dSP_958_p;
  wire       [31:0]   dSP_959_p;
  wire       [31:0]   dSP_960_p;
  wire       [31:0]   dSP_961_p;
  wire       [31:0]   dSP_962_p;
  wire       [31:0]   dSP_963_p;
  wire       [31:0]   dSP_964_p;
  wire       [31:0]   dSP_965_p;
  wire       [31:0]   dSP_966_p;
  wire       [31:0]   dSP_967_p;
  wire       [31:0]   dSP_968_p;
  wire       [31:0]   dSP_969_p;
  wire       [31:0]   dSP_970_p;
  wire       [31:0]   dSP_971_p;
  wire       [31:0]   dSP_972_p;
  wire       [31:0]   dSP_973_p;
  wire       [31:0]   dSP_974_p;
  wire       [31:0]   dSP_975_p;
  wire       [31:0]   dSP_976_p;
  wire       [31:0]   dSP_977_p;
  wire       [31:0]   dSP_978_p;
  wire       [31:0]   dSP_979_p;
  wire       [31:0]   dSP_980_p;
  wire       [31:0]   dSP_981_p;
  wire       [31:0]   dSP_982_p;
  wire       [31:0]   dSP_983_p;
  wire       [31:0]   dSP_984_p;
  wire       [31:0]   dSP_985_p;
  wire       [31:0]   dSP_986_p;
  wire       [31:0]   dSP_987_p;
  wire       [31:0]   dSP_988_p;
  wire       [31:0]   dSP_989_p;
  wire       [31:0]   dSP_990_p;
  wire       [31:0]   dSP_991_p;
  wire       [31:0]   dSP_992_p;
  wire       [31:0]   dSP_993_p;
  wire       [31:0]   dSP_994_p;
  wire       [31:0]   dSP_995_p;
  wire       [31:0]   dSP_996_p;
  wire       [31:0]   dSP_997_p;
  wire       [31:0]   dSP_998_p;
  wire       [31:0]   dSP_999_p;
  wire       [31:0]   dSP_1000_p;
  wire       [31:0]   dSP_1001_p;
  wire       [31:0]   dSP_1002_p;
  wire       [31:0]   dSP_1003_p;
  wire       [31:0]   dSP_1004_p;
  wire       [31:0]   dSP_1005_p;
  wire       [31:0]   dSP_1006_p;
  wire       [31:0]   dSP_1007_p;
  wire       [31:0]   dSP_1008_p;
  wire       [31:0]   dSP_1009_p;
  wire       [31:0]   dSP_1010_p;
  wire       [31:0]   dSP_1011_p;
  wire       [31:0]   dSP_1012_p;
  wire       [31:0]   dSP_1013_p;
  wire       [31:0]   dSP_1014_p;
  wire       [31:0]   dSP_1015_p;
  wire       [31:0]   dSP_1016_p;
  wire       [31:0]   dSP_1017_p;
  wire       [31:0]   dSP_1018_p;
  wire       [31:0]   dSP_1019_p;
  wire       [31:0]   dSP_1020_p;
  wire       [31:0]   dSP_1021_p;
  wire       [31:0]   dSP_1022_p;
  wire       [31:0]   dSP_1023_p;
  wire       [31:0]   dSP_1024_p;
  wire       [31:0]   dSP_1025_p;
  wire       [31:0]   dSP_1026_p;
  wire       [31:0]   dSP_1027_p;
  wire       [31:0]   dSP_1028_p;
  wire       [31:0]   dSP_1029_p;
  wire       [31:0]   dSP_1030_p;
  wire       [31:0]   dSP_1031_p;
  wire       [31:0]   dSP_1032_p;
  wire       [31:0]   dSP_1033_p;
  wire       [31:0]   dSP_1034_p;
  wire       [31:0]   dSP_1035_p;
  wire       [31:0]   dSP_1036_p;
  wire       [31:0]   dSP_1037_p;
  wire       [31:0]   dSP_1038_p;
  wire       [31:0]   dSP_1039_p;
  wire       [31:0]   dSP_1040_p;
  wire       [31:0]   dSP_1041_p;
  wire       [31:0]   dSP_1042_p;
  wire       [31:0]   dSP_1043_p;
  wire       [31:0]   dSP_1044_p;
  wire       [31:0]   dSP_1045_p;
  wire       [31:0]   dSP_1046_p;
  wire       [31:0]   dSP_1047_p;
  wire       [31:0]   dSP_1048_p;
  wire       [31:0]   dSP_1049_p;
  wire       [31:0]   dSP_1050_p;
  wire       [31:0]   dSP_1051_p;
  wire       [31:0]   dSP_1052_p;
  wire       [31:0]   dSP_1053_p;
  wire       [31:0]   dSP_1054_p;
  wire       [31:0]   dSP_1055_p;
  wire       [31:0]   dSP_1056_p;
  wire       [31:0]   dSP_1057_p;
  wire       [31:0]   dSP_1058_p;
  wire       [31:0]   dSP_1059_p;
  wire       [31:0]   dSP_1060_p;
  wire       [31:0]   dSP_1061_p;
  wire       [31:0]   dSP_1062_p;
  wire       [31:0]   dSP_1063_p;
  wire       [31:0]   dSP_1064_p;
  wire       [31:0]   dSP_1065_p;
  wire       [31:0]   dSP_1066_p;
  wire       [31:0]   dSP_1067_p;
  wire       [31:0]   dSP_1068_p;
  wire       [31:0]   dSP_1069_p;
  wire       [31:0]   dSP_1070_p;
  wire       [31:0]   dSP_1071_p;
  wire       [31:0]   dSP_1072_p;
  wire       [31:0]   dSP_1073_p;
  wire       [31:0]   dSP_1074_p;
  wire       [31:0]   dSP_1075_p;
  wire       [31:0]   dSP_1076_p;
  wire       [31:0]   dSP_1077_p;
  wire       [31:0]   dSP_1078_p;
  wire       [31:0]   dSP_1079_p;
  wire       [31:0]   dSP_1080_p;
  wire       [31:0]   dSP_1081_p;
  wire       [31:0]   dSP_1082_p;
  wire       [31:0]   dSP_1083_p;
  wire       [31:0]   dSP_1084_p;
  wire       [31:0]   dSP_1085_p;
  wire       [31:0]   dSP_1086_p;
  wire       [31:0]   dSP_1087_p;
  wire       [31:0]   dSP_1088_p;
  wire       [31:0]   dSP_1089_p;
  wire       [31:0]   dSP_1090_p;
  wire       [31:0]   dSP_1091_p;
  wire       [31:0]   dSP_1092_p;
  wire       [31:0]   dSP_1093_p;
  wire       [31:0]   dSP_1094_p;
  wire       [31:0]   dSP_1095_p;
  wire       [31:0]   dSP_1096_p;
  wire       [31:0]   dSP_1097_p;
  wire       [31:0]   dSP_1098_p;
  wire       [31:0]   dSP_1099_p;
  wire       [31:0]   dSP_1100_p;
  wire       [31:0]   dSP_1101_p;
  wire       [31:0]   dSP_1102_p;
  wire       [31:0]   dSP_1103_p;
  wire       [31:0]   dSP_1104_p;
  wire       [31:0]   dSP_1105_p;
  wire       [31:0]   dSP_1106_p;
  wire       [31:0]   dSP_1107_p;
  wire       [31:0]   dSP_1108_p;
  wire       [31:0]   dSP_1109_p;
  wire       [31:0]   dSP_1110_p;
  wire       [31:0]   dSP_1111_p;
  wire       [31:0]   dSP_1112_p;
  wire       [31:0]   dSP_1113_p;
  wire       [31:0]   dSP_1114_p;
  wire       [31:0]   dSP_1115_p;
  wire       [31:0]   dSP_1116_p;
  wire       [31:0]   dSP_1117_p;
  wire       [31:0]   dSP_1118_p;
  wire       [31:0]   dSP_1119_p;
  wire       [31:0]   dSP_1120_p;
  wire       [31:0]   dSP_1121_p;
  wire       [31:0]   dSP_1122_p;
  wire       [31:0]   dSP_1123_p;
  wire       [31:0]   dSP_1124_p;
  wire       [31:0]   dSP_1125_p;
  wire       [31:0]   dSP_1126_p;
  wire       [31:0]   dSP_1127_p;
  wire       [31:0]   dSP_1128_p;
  wire       [31:0]   dSP_1129_p;
  wire       [31:0]   dSP_1130_p;
  wire       [31:0]   dSP_1131_p;
  wire       [31:0]   dSP_1132_p;
  wire       [31:0]   dSP_1133_p;
  wire       [31:0]   dSP_1134_p;
  wire       [31:0]   dSP_1135_p;
  wire       [31:0]   dSP_1136_p;
  wire       [31:0]   dSP_1137_p;
  wire       [31:0]   dSP_1138_p;
  wire       [31:0]   dSP_1139_p;
  wire       [31:0]   dSP_1140_p;
  wire       [31:0]   dSP_1141_p;
  wire       [31:0]   dSP_1142_p;
  wire       [31:0]   dSP_1143_p;
  wire       [31:0]   dSP_1144_p;
  wire       [31:0]   dSP_1145_p;
  wire       [31:0]   dSP_1146_p;
  wire       [31:0]   dSP_1147_p;
  wire       [31:0]   dSP_1148_p;
  wire       [31:0]   dSP_1149_p;
  wire       [31:0]   dSP_1150_p;
  wire       [31:0]   dSP_1151_p;
  wire       [31:0]   dSP_1152_p;
  wire       [39:0]   addKernel_S;
  wire       [39:0]   addKernel_1_S;
  wire       [39:0]   addKernel_2_S;
  wire       [39:0]   addKernel_3_S;
  wire       [39:0]   addKernel_4_S;
  wire       [39:0]   addKernel_5_S;
  wire       [39:0]   addKernel_6_S;
  wire       [39:0]   addKernel_7_S;
  wire       [39:0]   addKernel_8_S;
  wire       [39:0]   addKernel_9_S;
  wire       [39:0]   addKernel_10_S;
  wire       [39:0]   addKernel_11_S;
  wire       [39:0]   addKernel_12_S;
  wire       [39:0]   addKernel_13_S;
  wire       [39:0]   addKernel_14_S;
  wire       [39:0]   addKernel_15_S;
  wire       [39:0]   addKernel_16_S;
  wire       [39:0]   addKernel_17_S;
  wire       [39:0]   addKernel_18_S;
  wire       [39:0]   addKernel_19_S;
  wire       [39:0]   addKernel_20_S;
  wire       [39:0]   addKernel_21_S;
  wire       [39:0]   addKernel_22_S;
  wire       [39:0]   addKernel_23_S;
  wire       [39:0]   addKernel_24_S;
  wire       [39:0]   addKernel_25_S;
  wire       [39:0]   addKernel_26_S;
  wire       [39:0]   addKernel_27_S;
  wire       [39:0]   addKernel_28_S;
  wire       [39:0]   addKernel_29_S;
  wire       [39:0]   addKernel_30_S;
  wire       [39:0]   addKernel_31_S;
  wire       [39:0]   addKernel_32_S;
  wire       [39:0]   addKernel_33_S;
  wire       [39:0]   addKernel_34_S;
  wire       [39:0]   addKernel_35_S;
  wire       [39:0]   addKernel_36_S;
  wire       [39:0]   addKernel_37_S;
  wire       [39:0]   addKernel_38_S;
  wire       [39:0]   addKernel_39_S;
  wire       [39:0]   addKernel_40_S;
  wire       [39:0]   addKernel_41_S;
  wire       [39:0]   addKernel_42_S;
  wire       [39:0]   addKernel_43_S;
  wire       [39:0]   addKernel_44_S;
  wire       [39:0]   addKernel_45_S;
  wire       [39:0]   addKernel_46_S;
  wire       [39:0]   addKernel_47_S;
  wire       [39:0]   addKernel_48_S;
  wire       [39:0]   addKernel_49_S;
  wire       [39:0]   addKernel_50_S;
  wire       [39:0]   addKernel_51_S;
  wire       [39:0]   addKernel_52_S;
  wire       [39:0]   addKernel_53_S;
  wire       [39:0]   addKernel_54_S;
  wire       [39:0]   addKernel_55_S;
  wire       [39:0]   addKernel_56_S;
  wire       [39:0]   addKernel_57_S;
  wire       [39:0]   addKernel_58_S;
  wire       [39:0]   addKernel_59_S;
  wire       [39:0]   addKernel_60_S;
  wire       [39:0]   addKernel_61_S;
  wire       [39:0]   addKernel_62_S;
  wire       [39:0]   addKernel_63_S;
  wire       [39:0]   addKernel_64_S;
  wire       [39:0]   addKernel_65_S;
  wire       [39:0]   addKernel_66_S;
  wire       [39:0]   addKernel_67_S;
  wire       [39:0]   addKernel_68_S;
  wire       [39:0]   addKernel_69_S;
  wire       [39:0]   addKernel_70_S;
  wire       [39:0]   addKernel_71_S;
  wire       [39:0]   addKernel_72_S;
  wire       [39:0]   addKernel_73_S;
  wire       [39:0]   addKernel_74_S;
  wire       [39:0]   addKernel_75_S;
  wire       [39:0]   addKernel_76_S;
  wire       [39:0]   addKernel_77_S;
  wire       [39:0]   addKernel_78_S;
  wire       [39:0]   addKernel_79_S;
  wire       [39:0]   addKernel_80_S;
  wire       [39:0]   addKernel_81_S;
  wire       [39:0]   addKernel_82_S;
  wire       [39:0]   addKernel_83_S;
  wire       [39:0]   addKernel_84_S;
  wire       [39:0]   addKernel_85_S;
  wire       [39:0]   addKernel_86_S;
  wire       [39:0]   addKernel_87_S;
  wire       [39:0]   addKernel_88_S;
  wire       [39:0]   addKernel_89_S;
  wire       [39:0]   addKernel_90_S;
  wire       [39:0]   addKernel_91_S;
  wire       [39:0]   addKernel_92_S;
  wire       [39:0]   addKernel_93_S;
  wire       [39:0]   addKernel_94_S;
  wire       [39:0]   addKernel_95_S;
  wire       [39:0]   addKernel_96_S;
  wire       [39:0]   addKernel_97_S;
  wire       [39:0]   addKernel_98_S;
  wire       [39:0]   addKernel_99_S;
  wire       [39:0]   addKernel_100_S;
  wire       [39:0]   addKernel_101_S;
  wire       [39:0]   addKernel_102_S;
  wire       [39:0]   addKernel_103_S;
  wire       [39:0]   addKernel_104_S;
  wire       [39:0]   addKernel_105_S;
  wire       [39:0]   addKernel_106_S;
  wire       [39:0]   addKernel_107_S;
  wire       [39:0]   addKernel_108_S;
  wire       [39:0]   addKernel_109_S;
  wire       [39:0]   addKernel_110_S;
  wire       [39:0]   addKernel_111_S;
  wire       [39:0]   addKernel_112_S;
  wire       [39:0]   addKernel_113_S;
  wire       [39:0]   addKernel_114_S;
  wire       [39:0]   addKernel_115_S;
  wire       [39:0]   addKernel_116_S;
  wire       [39:0]   addKernel_117_S;
  wire       [39:0]   addKernel_118_S;
  wire       [39:0]   addKernel_119_S;
  wire       [39:0]   addKernel_120_S;
  wire       [39:0]   addKernel_121_S;
  wire       [39:0]   addKernel_122_S;
  wire       [39:0]   addKernel_123_S;
  wire       [39:0]   addKernel_124_S;
  wire       [39:0]   addKernel_125_S;
  wire       [39:0]   addKernel_126_S;
  wire       [39:0]   addKernel_127_S;
  wire       [47:0]   xAddTimes_136_S;
  wire       [47:0]   xAddTimes_137_S;
  wire       [47:0]   xAddTimes_138_S;
  wire       [47:0]   xAddTimes_139_S;
  wire       [47:0]   xAddTimes_140_S;
  wire       [47:0]   xAddTimes_141_S;
  wire       [47:0]   xAddTimes_142_S;
  wire       [47:0]   xAddTimes_143_S;
  wire       [31:0]   xAddChannelTimes_16_S;
  wire       [31:0]   xAddChannelTimes_17_S;
  wire       [31:0]   xAddChannelTimes_18_S;
  wire       [31:0]   xAddChannelTimes_19_S;
  wire       [31:0]   xAddChannelTimes_20_S;
  wire       [31:0]   xAddChannelTimes_21_S;
  wire       [31:0]   xAddChannelTimes_22_S;
  wire       [31:0]   xAddChannelTimes_23_S;
  wire       [31:0]   xAddChannelTimes_24_S;
  wire       [31:0]   xAddChannelTimes_25_S;
  wire       [31:0]   xAddChannelTimes_26_S;
  wire       [31:0]   xAddChannelTimes_27_S;
  wire       [31:0]   xAddChannelTimes_28_S;
  wire       [31:0]   xAddChannelTimes_29_S;
  wire       [31:0]   xAddChannelTimes_30_S;
  wire       [31:0]   xAddChannelTimes_31_S;
  wire       [127:0]  quan_1_dataOut;
  wire                stride_1_sData_ready;
  wire                stride_1_mData_valid;
  wire       [127:0]  stride_1_mData_payload;
  wire                stride_1_sReady;
  wire                stride_1_complete;
  wire                stride_1_last;
  wire       [127:0]  _zz__zz_1_port;
  wire                _zz__zz_1_port_1;
  wire                _zz__zz_b_9;
  wire       [127:0]  _zz__zz_2_port;
  wire                _zz__zz_2_port_1;
  wire                _zz__zz_b_19;
  wire       [127:0]  _zz__zz_3_port;
  wire                _zz__zz_3_port_1;
  wire                _zz__zz_b_29;
  wire       [127:0]  _zz__zz_4_port;
  wire                _zz__zz_4_port_1;
  wire                _zz__zz_b_39;
  wire       [127:0]  _zz__zz_5_port;
  wire                _zz__zz_5_port_1;
  wire                _zz__zz_b_49;
  wire       [127:0]  _zz__zz_6_port;
  wire                _zz__zz_6_port_1;
  wire                _zz__zz_b_59;
  wire       [127:0]  _zz__zz_7_port;
  wire                _zz__zz_7_port_1;
  wire                _zz__zz_b_69;
  wire       [127:0]  _zz__zz_8_port;
  wire                _zz__zz_8_port_1;
  wire                _zz__zz_b_79;
  wire       [127:0]  _zz__zz_9_port;
  wire                _zz__zz_9_port_1;
  wire                _zz__zz_b_89;
  reg        [1:0]    _zz_convType;
  wire       [127:0]  _zz_b;
  wire       [127:0]  _zz_b_1;
  wire       [127:0]  _zz_b_2;
  wire       [127:0]  _zz_b_3;
  wire       [127:0]  _zz_b_4;
  wire       [127:0]  _zz_b_5;
  wire       [127:0]  _zz_b_6;
  wire       [127:0]  _zz_b_7;
  wire       [127:0]  _zz_b_8;
  reg        [127:0]  _zz_b_9;
  reg        [127:0]  _zz_b_10;
  reg        [127:0]  _zz_b_11;
  reg        [127:0]  _zz_b_12;
  reg        [127:0]  _zz_b_13;
  reg        [127:0]  _zz_b_14;
  reg        [127:0]  _zz_b_15;
  reg        [127:0]  _zz_b_16;
  reg        [127:0]  _zz_b_17;
  reg        [127:0]  _zz_b_18;
  reg        [127:0]  _zz_b_19;
  reg        [127:0]  _zz_b_20;
  reg        [127:0]  _zz_b_21;
  reg        [127:0]  _zz_b_22;
  reg        [127:0]  _zz_b_23;
  reg        [127:0]  _zz_b_24;
  reg        [127:0]  _zz_b_25;
  reg        [127:0]  _zz_b_26;
  reg        [127:0]  _zz_b_27;
  reg        [127:0]  _zz_b_28;
  reg        [127:0]  _zz_b_29;
  reg        [127:0]  _zz_b_30;
  reg        [127:0]  _zz_b_31;
  reg        [127:0]  _zz_b_32;
  reg        [127:0]  _zz_b_33;
  reg        [127:0]  _zz_b_34;
  reg        [127:0]  _zz_b_35;
  reg        [127:0]  _zz_b_36;
  reg        [127:0]  _zz_b_37;
  reg        [127:0]  _zz_b_38;
  reg        [127:0]  _zz_b_39;
  reg        [127:0]  _zz_b_40;
  reg        [127:0]  _zz_b_41;
  reg        [127:0]  _zz_b_42;
  reg        [127:0]  _zz_b_43;
  reg        [127:0]  _zz_b_44;
  reg        [127:0]  _zz_b_45;
  reg        [127:0]  _zz_b_46;
  reg        [127:0]  _zz_b_47;
  reg        [127:0]  _zz_b_48;
  reg        [127:0]  _zz_b_49;
  reg        [127:0]  _zz_b_50;
  reg        [127:0]  _zz_b_51;
  reg        [127:0]  _zz_b_52;
  reg        [127:0]  _zz_b_53;
  reg        [127:0]  _zz_b_54;
  reg        [127:0]  _zz_b_55;
  reg        [127:0]  _zz_b_56;
  reg        [127:0]  _zz_b_57;
  reg        [127:0]  _zz_b_58;
  reg        [127:0]  _zz_b_59;
  reg        [127:0]  _zz_b_60;
  reg        [127:0]  _zz_b_61;
  reg        [127:0]  _zz_b_62;
  reg        [127:0]  _zz_b_63;
  reg        [127:0]  _zz_b_64;
  reg        [127:0]  _zz_b_65;
  reg        [127:0]  _zz_b_66;
  reg        [127:0]  _zz_b_67;
  reg        [127:0]  _zz_b_68;
  reg        [127:0]  _zz_b_69;
  reg        [127:0]  _zz_b_70;
  reg        [127:0]  _zz_b_71;
  reg        [127:0]  _zz_b_72;
  reg        [127:0]  _zz_b_73;
  reg        [127:0]  _zz_b_74;
  reg        [127:0]  _zz_b_75;
  reg        [127:0]  _zz_b_76;
  reg        [127:0]  _zz_b_77;
  reg        [127:0]  _zz_b_78;
  reg        [127:0]  _zz_b_79;
  reg        [127:0]  _zz_b_80;
  reg        [127:0]  _zz_b_81;
  reg        [127:0]  _zz_b_82;
  reg        [127:0]  _zz_b_83;
  reg        [127:0]  _zz_b_84;
  reg        [127:0]  _zz_b_85;
  reg        [127:0]  _zz_b_86;
  reg        [127:0]  _zz_b_87;
  reg        [127:0]  _zz_b_88;
  reg        [127:0]  _zz_b_89;
  reg        [127:0]  _zz_b_90;
  reg        [127:0]  _zz_b_91;
  reg        [127:0]  _zz_b_92;
  reg        [127:0]  _zz_b_93;
  reg        [127:0]  _zz_b_94;
  reg        [127:0]  _zz_b_95;
  reg        [127:0]  _zz_b_96;
  reg        [127:0]  _zz_b_97;
  reg        [127:0]  _zz_b_98;
  wire       [47:0]   _zz_A;
  wire       [47:0]   _zz_A_1;
  wire       [47:0]   _zz_A_2;
  wire       [47:0]   _zz_A_3;
  wire       [47:0]   _zz_A_4;
  wire       [47:0]   _zz_A_5;
  wire       [47:0]   _zz_A_6;
  wire       [47:0]   _zz_A_7;
  (* ram_style = "block" *) reg [127:0] _zz_1 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_2 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_3 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_4 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_5 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_6 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_7 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_8 [0:31];
  (* ram_style = "block" *) reg [127:0] _zz_9 [0:31];

  assign _zz__zz_1_port = waXpmSyncFifo_9_dout;
  assign _zz__zz_b_9 = 1'b1;
  assign _zz__zz_2_port = waXpmSyncFifo_10_dout;
  assign _zz__zz_b_19 = 1'b1;
  assign _zz__zz_3_port = waXpmSyncFifo_11_dout;
  assign _zz__zz_b_29 = 1'b1;
  assign _zz__zz_4_port = waXpmSyncFifo_12_dout;
  assign _zz__zz_b_39 = 1'b1;
  assign _zz__zz_5_port = waXpmSyncFifo_13_dout;
  assign _zz__zz_b_49 = 1'b1;
  assign _zz__zz_6_port = waXpmSyncFifo_14_dout;
  assign _zz__zz_b_59 = 1'b1;
  assign _zz__zz_7_port = waXpmSyncFifo_15_dout;
  assign _zz__zz_b_69 = 1'b1;
  assign _zz__zz_8_port = waXpmSyncFifo_16_dout;
  assign _zz__zz_b_79 = 1'b1;
  assign _zz__zz_9_port = waXpmSyncFifo_17_dout;
  assign _zz__zz_b_89 = 1'b1;
  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_1[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_1_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_9) begin
      _zz__zz_1_port1 <= _zz_1[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_2[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_2_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_19) begin
      _zz__zz_2_port1 <= _zz_2[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_3[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_3_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_29) begin
      _zz__zz_3_port1 <= _zz_3[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_4[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_4_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_39) begin
      _zz__zz_4_port1 <= _zz_4[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_5[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_5_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_49) begin
      _zz__zz_5_port1 <= _zz_5[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_6[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_6_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_59) begin
      _zz__zz_6_port1 <= _zz_6[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_7[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_7_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_69) begin
      _zz__zz_7_port1 <= _zz_7[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_8[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_8_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_79) begin
      _zz__zz_8_port1 <= _zz_8[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  always @(posedge clk) begin
    if(convComputeCtrl_1_featureMemWriteReady) begin
      _zz_9[convComputeCtrl_1_featureMemWriteAddr] <= _zz__zz_9_port;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_b_89) begin
      _zz__zz_9_port1 <= _zz_9[convComputeCtrl_1_featureMemReadAddr];
    end
  end

  ChannelIncr channelIncr_1 (
    .sData_valid   (sFeatureFirstLayerData_valid       ), //i
    .sData_ready   (channelIncr_1_sData_ready          ), //o
    .sData_payload (sFeatureFirstLayerData_payload[7:0]), //i
    .mData_valid   (channelIncr_1_mData_valid          ), //o
    .mData_ready   (channelIncr_1_mData_ready          ), //i
    .mData_payload (channelIncr_1_mData_payload[127:0] )  //o
  );
  DataGenerate dataGenerate_1 (
    .sData_valid           (dataGenerate_1_sData_valid                 ), //i
    .sData_ready           (dataGenerate_1_sData_ready                 ), //o
    .sData_payload         (dataGenerate_1_sData_payload[127:0]        ), //i
    .start                 (startCu                                    ), //i
    .enPadding             (enPadding                                  ), //i
    .channelIn             (channelIn[11:0]                            ), //i
    .rowNumIn              (rowNumIn[9:0]                              ), //i
    .colNumIn              (colNumIn[9:0]                              ), //i
    .zeroDara              (zeroDara[7:0]                              ), //i
    .zeroNum               (zeroNum                                    ), //i
    .mData_mData_0_valid   (dataGenerate_1_mData_mData_0_valid         ), //o
    .mData_mData_0_payload (dataGenerate_1_mData_mData_0_payload[127:0]), //o
    .mData_mData_1_valid   (dataGenerate_1_mData_mData_1_valid         ), //o
    .mData_mData_1_payload (dataGenerate_1_mData_mData_1_payload[127:0]), //o
    .mData_mData_2_valid   (dataGenerate_1_mData_mData_2_valid         ), //o
    .mData_mData_2_payload (dataGenerate_1_mData_mData_2_payload[127:0]), //o
    .mData_mData_3_valid   (dataGenerate_1_mData_mData_3_valid         ), //o
    .mData_mData_3_payload (dataGenerate_1_mData_mData_3_payload[127:0]), //o
    .mData_mData_4_valid   (dataGenerate_1_mData_mData_4_valid         ), //o
    .mData_mData_4_payload (dataGenerate_1_mData_mData_4_payload[127:0]), //o
    .mData_mData_5_valid   (dataGenerate_1_mData_mData_5_valid         ), //o
    .mData_mData_5_payload (dataGenerate_1_mData_mData_5_payload[127:0]), //o
    .mData_mData_6_valid   (dataGenerate_1_mData_mData_6_valid         ), //o
    .mData_mData_6_payload (dataGenerate_1_mData_mData_6_payload[127:0]), //o
    .mData_mData_7_valid   (dataGenerate_1_mData_mData_7_valid         ), //o
    .mData_mData_7_payload (dataGenerate_1_mData_mData_7_payload[127:0]), //o
    .mData_mData_8_valid   (dataGenerate_1_mData_mData_8_valid         ), //o
    .mData_mData_8_payload (dataGenerate_1_mData_mData_8_payload[127:0]), //o
    .mData_ready           (waXpmSyncFifo_9_sReady                     ), //i
    .convType              (_zz_convType[1:0]                          ), //i
    .reset                 (reset                                      ), //i
    .clk                   (clk                                        ), //i
    .softReset             (softReset                                  )  //i
  );
  ConvComputeCtrl convComputeCtrl_1 (
    .start                (startCu                                   ), //i
    .mDataValid           (convComputeCtrl_1_mDataValid              ), //o
    .mDataReady           (stride_1_sReady                           ), //i
    .normPreValid         (convComputeCtrl_1_normPreValid            ), //o
    .sDataReady           (waXpmSyncFifo_9_mReady                    ), //i
    .rowNumIn             (rowNumIn[9:0]                             ), //i
    .colNumIn             (colNumIn[9:0]                             ), //i
    .channelIn            (channelIn[11:0]                           ), //i
    .channelOut           (channelOut[11:0]                          ), //i
    .featureMemReadAddr   (convComputeCtrl_1_featureMemReadAddr[4:0] ), //o
    .featureMemWriteAddr  (convComputeCtrl_1_featureMemWriteAddr[4:0]), //o
    .featureMemWriteReady (convComputeCtrl_1_featureMemWriteReady    ), //o
    .weightReadAddr_0     (convComputeCtrl_1_weightReadAddr_0[8:0]   ), //o
    .weightReadAddr_1     (convComputeCtrl_1_weightReadAddr_1[8:0]   ), //o
    .weightReadAddr_2     (convComputeCtrl_1_weightReadAddr_2[8:0]   ), //o
    .weightReadAddr_3     (convComputeCtrl_1_weightReadAddr_3[8:0]   ), //o
    .weightReadAddr_4     (convComputeCtrl_1_weightReadAddr_4[8:0]   ), //o
    .weightReadAddr_5     (convComputeCtrl_1_weightReadAddr_5[8:0]   ), //o
    .weightReadAddr_6     (convComputeCtrl_1_weightReadAddr_6[8:0]   ), //o
    .weightReadAddr_7     (convComputeCtrl_1_weightReadAddr_7[8:0]   ), //o
    .weightReadAddr_8     (convComputeCtrl_1_weightReadAddr_8[8:0]   ), //o
    .biasReadAddr         (convComputeCtrl_1_biasReadAddr[5:0]       ), //o
    .scaleReadAddr        (convComputeCtrl_1_scaleReadAddr[5:0]      ), //o
    .shiftReadAddr        (convComputeCtrl_1_shiftReadAddr[5:0]      ), //o
    .activationEn         (enActivation                              ), //i
    .sCount               (convComputeCtrl_1_sCount[12:0]            ), //o
    .mCount               (convComputeCtrl_1_mCount[12:0]            ), //o
    .convType             (_zz_convType[1:0]                         ), //i
    .clk                  (clk                                       ), //i
    .reset                (reset                                     ), //i
    .softReset            (softReset                                 )  //i
  );
  LoadWeight loadWeight_1 (
    .start             (startPa                                ), //i
    .sData_valid       (sParaData_valid                        ), //i
    .sData_ready       (loadWeight_1_sData_ready               ), //o
    .sData_payload     (sParaData_payload[127:0]               ), //i
    .weightNum         (weightNum[12:0]                        ), //i
    .quanNum           (quanNum[7:0]                           ), //i
    .weightRead_0_addr (convComputeCtrl_1_weightReadAddr_0[8:0]), //i
    .weightRead_0_data (loadWeight_1_weightRead_0_data[2047:0] ), //o
    .weightRead_1_addr (convComputeCtrl_1_weightReadAddr_1[8:0]), //i
    .weightRead_1_data (loadWeight_1_weightRead_1_data[2047:0] ), //o
    .weightRead_2_addr (convComputeCtrl_1_weightReadAddr_2[8:0]), //i
    .weightRead_2_data (loadWeight_1_weightRead_2_data[2047:0] ), //o
    .weightRead_3_addr (convComputeCtrl_1_weightReadAddr_3[8:0]), //i
    .weightRead_3_data (loadWeight_1_weightRead_3_data[2047:0] ), //o
    .weightRead_4_addr (convComputeCtrl_1_weightReadAddr_4[8:0]), //i
    .weightRead_4_data (loadWeight_1_weightRead_4_data[2047:0] ), //o
    .weightRead_5_addr (convComputeCtrl_1_weightReadAddr_5[8:0]), //i
    .weightRead_5_data (loadWeight_1_weightRead_5_data[2047:0] ), //o
    .weightRead_6_addr (convComputeCtrl_1_weightReadAddr_6[8:0]), //i
    .weightRead_6_data (loadWeight_1_weightRead_6_data[2047:0] ), //o
    .weightRead_7_addr (convComputeCtrl_1_weightReadAddr_7[8:0]), //i
    .weightRead_7_data (loadWeight_1_weightRead_7_data[2047:0] ), //o
    .weightRead_8_addr (convComputeCtrl_1_weightReadAddr_8[8:0]), //i
    .weightRead_8_data (loadWeight_1_weightRead_8_data[2047:0] ), //o
    .biasRead_addr     (convComputeCtrl_1_biasReadAddr[5:0]    ), //i
    .biasRead_data     (loadWeight_1_biasRead_data[511:0]      ), //o
    .scaleRead_addr    (convComputeCtrl_1_scaleReadAddr[5:0]   ), //i
    .scaleRead_data    (loadWeight_1_scaleRead_data[511:0]     ), //o
    .shiftRead_addr    (convComputeCtrl_1_shiftReadAddr[5:0]   ), //i
    .shiftRead_data    (loadWeight_1_shiftRead_data[511:0]     ), //o
    .copyWeightDone    (loadWeight_1_copyWeightDone            ), //o
    .convType          (convType[1:0]                          ), //i
    .channelIn         (channelIn[11:0]                        ), //i
    .channelOut        (channelOut[11:0]                       ), //i
    .clk               (clk                                    ), //i
    .reset             (reset                                  ), //i
    .softReset         (softReset                              )  //i
  );
  WaXpmSyncFifo waXpmSyncFifo_9 (
    .sCount         (waXpmSyncFifo_9_sCount[13:0]               ), //i
    .mCount         (waXpmSyncFifo_9_mCount[13:0]               ), //i
    .sReady         (waXpmSyncFifo_9_sReady                     ), //o
    .mReady         (waXpmSyncFifo_9_mReady                     ), //o
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_0_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_0_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_9_dout[127:0]                ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_10 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_1_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_1_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_10_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_11 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_2_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_2_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_11_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_12 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_3_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_3_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_12_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_13 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_4_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_4_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_13_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_14 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_5_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_5_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_14_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_15 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_6_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_6_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_15_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_16 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_7_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_7_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_16_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  WaXpmSyncFifo_1 waXpmSyncFifo_17 (
    .reset          (reset                                      ), //i
    .clk            (clk                                        ), //i
    .dataIn_valid   (dataGenerate_1_mData_mData_8_valid         ), //i
    .dataIn_payload (dataGenerate_1_mData_mData_8_payload[127:0]), //i
    .rd_en          (convComputeCtrl_1_featureMemWriteReady     ), //i
    .dout           (waXpmSyncFifo_17_dout[127:0]               ), //o
    .softReset      (softReset                                  )  //i
  );
  DSP dSP_1 (
    .a   (dSP_1_a[7:0] ), //i
    .d   (dSP_1_d[7:0] ), //i
    .b   (dSP_1_b[7:0] ), //i
    .p   (dSP_1_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_2 (
    .a   (dSP_2_a[7:0] ), //i
    .d   (dSP_2_d[7:0] ), //i
    .b   (dSP_2_b[7:0] ), //i
    .p   (dSP_2_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_3 (
    .a   (dSP_3_a[7:0] ), //i
    .d   (dSP_3_d[7:0] ), //i
    .b   (dSP_3_b[7:0] ), //i
    .p   (dSP_3_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_4 (
    .a   (dSP_4_a[7:0] ), //i
    .d   (dSP_4_d[7:0] ), //i
    .b   (dSP_4_b[7:0] ), //i
    .p   (dSP_4_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_5 (
    .a   (dSP_5_a[7:0] ), //i
    .d   (dSP_5_d[7:0] ), //i
    .b   (dSP_5_b[7:0] ), //i
    .p   (dSP_5_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_6 (
    .a   (dSP_6_a[7:0] ), //i
    .d   (dSP_6_d[7:0] ), //i
    .b   (dSP_6_b[7:0] ), //i
    .p   (dSP_6_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_7 (
    .a   (dSP_7_a[7:0] ), //i
    .d   (dSP_7_d[7:0] ), //i
    .b   (dSP_7_b[7:0] ), //i
    .p   (dSP_7_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_8 (
    .a   (dSP_8_a[7:0] ), //i
    .d   (dSP_8_d[7:0] ), //i
    .b   (dSP_8_b[7:0] ), //i
    .p   (dSP_8_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_9 (
    .a   (dSP_9_a[7:0] ), //i
    .d   (dSP_9_d[7:0] ), //i
    .b   (dSP_9_b[7:0] ), //i
    .p   (dSP_9_p[31:0]), //o
    .CLK (clk          )  //i
  );
  DSP dSP_10 (
    .a   (dSP_10_a[7:0] ), //i
    .d   (dSP_10_d[7:0] ), //i
    .b   (dSP_10_b[7:0] ), //i
    .p   (dSP_10_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_11 (
    .a   (dSP_11_a[7:0] ), //i
    .d   (dSP_11_d[7:0] ), //i
    .b   (dSP_11_b[7:0] ), //i
    .p   (dSP_11_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_12 (
    .a   (dSP_12_a[7:0] ), //i
    .d   (dSP_12_d[7:0] ), //i
    .b   (dSP_12_b[7:0] ), //i
    .p   (dSP_12_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_13 (
    .a   (dSP_13_a[7:0] ), //i
    .d   (dSP_13_d[7:0] ), //i
    .b   (dSP_13_b[7:0] ), //i
    .p   (dSP_13_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_14 (
    .a   (dSP_14_a[7:0] ), //i
    .d   (dSP_14_d[7:0] ), //i
    .b   (dSP_14_b[7:0] ), //i
    .p   (dSP_14_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_15 (
    .a   (dSP_15_a[7:0] ), //i
    .d   (dSP_15_d[7:0] ), //i
    .b   (dSP_15_b[7:0] ), //i
    .p   (dSP_15_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_16 (
    .a   (dSP_16_a[7:0] ), //i
    .d   (dSP_16_d[7:0] ), //i
    .b   (dSP_16_b[7:0] ), //i
    .p   (dSP_16_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_17 (
    .a   (dSP_17_a[7:0] ), //i
    .d   (dSP_17_d[7:0] ), //i
    .b   (dSP_17_b[7:0] ), //i
    .p   (dSP_17_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_18 (
    .a   (dSP_18_a[7:0] ), //i
    .d   (dSP_18_d[7:0] ), //i
    .b   (dSP_18_b[7:0] ), //i
    .p   (dSP_18_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_19 (
    .a   (dSP_19_a[7:0] ), //i
    .d   (dSP_19_d[7:0] ), //i
    .b   (dSP_19_b[7:0] ), //i
    .p   (dSP_19_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_20 (
    .a   (dSP_20_a[7:0] ), //i
    .d   (dSP_20_d[7:0] ), //i
    .b   (dSP_20_b[7:0] ), //i
    .p   (dSP_20_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_21 (
    .a   (dSP_21_a[7:0] ), //i
    .d   (dSP_21_d[7:0] ), //i
    .b   (dSP_21_b[7:0] ), //i
    .p   (dSP_21_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_22 (
    .a   (dSP_22_a[7:0] ), //i
    .d   (dSP_22_d[7:0] ), //i
    .b   (dSP_22_b[7:0] ), //i
    .p   (dSP_22_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_23 (
    .a   (dSP_23_a[7:0] ), //i
    .d   (dSP_23_d[7:0] ), //i
    .b   (dSP_23_b[7:0] ), //i
    .p   (dSP_23_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_24 (
    .a   (dSP_24_a[7:0] ), //i
    .d   (dSP_24_d[7:0] ), //i
    .b   (dSP_24_b[7:0] ), //i
    .p   (dSP_24_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_25 (
    .a   (dSP_25_a[7:0] ), //i
    .d   (dSP_25_d[7:0] ), //i
    .b   (dSP_25_b[7:0] ), //i
    .p   (dSP_25_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_26 (
    .a   (dSP_26_a[7:0] ), //i
    .d   (dSP_26_d[7:0] ), //i
    .b   (dSP_26_b[7:0] ), //i
    .p   (dSP_26_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_27 (
    .a   (dSP_27_a[7:0] ), //i
    .d   (dSP_27_d[7:0] ), //i
    .b   (dSP_27_b[7:0] ), //i
    .p   (dSP_27_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_28 (
    .a   (dSP_28_a[7:0] ), //i
    .d   (dSP_28_d[7:0] ), //i
    .b   (dSP_28_b[7:0] ), //i
    .p   (dSP_28_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_29 (
    .a   (dSP_29_a[7:0] ), //i
    .d   (dSP_29_d[7:0] ), //i
    .b   (dSP_29_b[7:0] ), //i
    .p   (dSP_29_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_30 (
    .a   (dSP_30_a[7:0] ), //i
    .d   (dSP_30_d[7:0] ), //i
    .b   (dSP_30_b[7:0] ), //i
    .p   (dSP_30_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_31 (
    .a   (dSP_31_a[7:0] ), //i
    .d   (dSP_31_d[7:0] ), //i
    .b   (dSP_31_b[7:0] ), //i
    .p   (dSP_31_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_32 (
    .a   (dSP_32_a[7:0] ), //i
    .d   (dSP_32_d[7:0] ), //i
    .b   (dSP_32_b[7:0] ), //i
    .p   (dSP_32_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_33 (
    .a   (dSP_33_a[7:0] ), //i
    .d   (dSP_33_d[7:0] ), //i
    .b   (dSP_33_b[7:0] ), //i
    .p   (dSP_33_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_34 (
    .a   (dSP_34_a[7:0] ), //i
    .d   (dSP_34_d[7:0] ), //i
    .b   (dSP_34_b[7:0] ), //i
    .p   (dSP_34_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_35 (
    .a   (dSP_35_a[7:0] ), //i
    .d   (dSP_35_d[7:0] ), //i
    .b   (dSP_35_b[7:0] ), //i
    .p   (dSP_35_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_36 (
    .a   (dSP_36_a[7:0] ), //i
    .d   (dSP_36_d[7:0] ), //i
    .b   (dSP_36_b[7:0] ), //i
    .p   (dSP_36_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_37 (
    .a   (dSP_37_a[7:0] ), //i
    .d   (dSP_37_d[7:0] ), //i
    .b   (dSP_37_b[7:0] ), //i
    .p   (dSP_37_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_38 (
    .a   (dSP_38_a[7:0] ), //i
    .d   (dSP_38_d[7:0] ), //i
    .b   (dSP_38_b[7:0] ), //i
    .p   (dSP_38_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_39 (
    .a   (dSP_39_a[7:0] ), //i
    .d   (dSP_39_d[7:0] ), //i
    .b   (dSP_39_b[7:0] ), //i
    .p   (dSP_39_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_40 (
    .a   (dSP_40_a[7:0] ), //i
    .d   (dSP_40_d[7:0] ), //i
    .b   (dSP_40_b[7:0] ), //i
    .p   (dSP_40_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_41 (
    .a   (dSP_41_a[7:0] ), //i
    .d   (dSP_41_d[7:0] ), //i
    .b   (dSP_41_b[7:0] ), //i
    .p   (dSP_41_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_42 (
    .a   (dSP_42_a[7:0] ), //i
    .d   (dSP_42_d[7:0] ), //i
    .b   (dSP_42_b[7:0] ), //i
    .p   (dSP_42_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_43 (
    .a   (dSP_43_a[7:0] ), //i
    .d   (dSP_43_d[7:0] ), //i
    .b   (dSP_43_b[7:0] ), //i
    .p   (dSP_43_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_44 (
    .a   (dSP_44_a[7:0] ), //i
    .d   (dSP_44_d[7:0] ), //i
    .b   (dSP_44_b[7:0] ), //i
    .p   (dSP_44_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_45 (
    .a   (dSP_45_a[7:0] ), //i
    .d   (dSP_45_d[7:0] ), //i
    .b   (dSP_45_b[7:0] ), //i
    .p   (dSP_45_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_46 (
    .a   (dSP_46_a[7:0] ), //i
    .d   (dSP_46_d[7:0] ), //i
    .b   (dSP_46_b[7:0] ), //i
    .p   (dSP_46_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_47 (
    .a   (dSP_47_a[7:0] ), //i
    .d   (dSP_47_d[7:0] ), //i
    .b   (dSP_47_b[7:0] ), //i
    .p   (dSP_47_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_48 (
    .a   (dSP_48_a[7:0] ), //i
    .d   (dSP_48_d[7:0] ), //i
    .b   (dSP_48_b[7:0] ), //i
    .p   (dSP_48_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_49 (
    .a   (dSP_49_a[7:0] ), //i
    .d   (dSP_49_d[7:0] ), //i
    .b   (dSP_49_b[7:0] ), //i
    .p   (dSP_49_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_50 (
    .a   (dSP_50_a[7:0] ), //i
    .d   (dSP_50_d[7:0] ), //i
    .b   (dSP_50_b[7:0] ), //i
    .p   (dSP_50_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_51 (
    .a   (dSP_51_a[7:0] ), //i
    .d   (dSP_51_d[7:0] ), //i
    .b   (dSP_51_b[7:0] ), //i
    .p   (dSP_51_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_52 (
    .a   (dSP_52_a[7:0] ), //i
    .d   (dSP_52_d[7:0] ), //i
    .b   (dSP_52_b[7:0] ), //i
    .p   (dSP_52_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_53 (
    .a   (dSP_53_a[7:0] ), //i
    .d   (dSP_53_d[7:0] ), //i
    .b   (dSP_53_b[7:0] ), //i
    .p   (dSP_53_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_54 (
    .a   (dSP_54_a[7:0] ), //i
    .d   (dSP_54_d[7:0] ), //i
    .b   (dSP_54_b[7:0] ), //i
    .p   (dSP_54_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_55 (
    .a   (dSP_55_a[7:0] ), //i
    .d   (dSP_55_d[7:0] ), //i
    .b   (dSP_55_b[7:0] ), //i
    .p   (dSP_55_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_56 (
    .a   (dSP_56_a[7:0] ), //i
    .d   (dSP_56_d[7:0] ), //i
    .b   (dSP_56_b[7:0] ), //i
    .p   (dSP_56_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_57 (
    .a   (dSP_57_a[7:0] ), //i
    .d   (dSP_57_d[7:0] ), //i
    .b   (dSP_57_b[7:0] ), //i
    .p   (dSP_57_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_58 (
    .a   (dSP_58_a[7:0] ), //i
    .d   (dSP_58_d[7:0] ), //i
    .b   (dSP_58_b[7:0] ), //i
    .p   (dSP_58_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_59 (
    .a   (dSP_59_a[7:0] ), //i
    .d   (dSP_59_d[7:0] ), //i
    .b   (dSP_59_b[7:0] ), //i
    .p   (dSP_59_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_60 (
    .a   (dSP_60_a[7:0] ), //i
    .d   (dSP_60_d[7:0] ), //i
    .b   (dSP_60_b[7:0] ), //i
    .p   (dSP_60_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_61 (
    .a   (dSP_61_a[7:0] ), //i
    .d   (dSP_61_d[7:0] ), //i
    .b   (dSP_61_b[7:0] ), //i
    .p   (dSP_61_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_62 (
    .a   (dSP_62_a[7:0] ), //i
    .d   (dSP_62_d[7:0] ), //i
    .b   (dSP_62_b[7:0] ), //i
    .p   (dSP_62_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_63 (
    .a   (dSP_63_a[7:0] ), //i
    .d   (dSP_63_d[7:0] ), //i
    .b   (dSP_63_b[7:0] ), //i
    .p   (dSP_63_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_64 (
    .a   (dSP_64_a[7:0] ), //i
    .d   (dSP_64_d[7:0] ), //i
    .b   (dSP_64_b[7:0] ), //i
    .p   (dSP_64_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_65 (
    .a   (dSP_65_a[7:0] ), //i
    .d   (dSP_65_d[7:0] ), //i
    .b   (dSP_65_b[7:0] ), //i
    .p   (dSP_65_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_66 (
    .a   (dSP_66_a[7:0] ), //i
    .d   (dSP_66_d[7:0] ), //i
    .b   (dSP_66_b[7:0] ), //i
    .p   (dSP_66_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_67 (
    .a   (dSP_67_a[7:0] ), //i
    .d   (dSP_67_d[7:0] ), //i
    .b   (dSP_67_b[7:0] ), //i
    .p   (dSP_67_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_68 (
    .a   (dSP_68_a[7:0] ), //i
    .d   (dSP_68_d[7:0] ), //i
    .b   (dSP_68_b[7:0] ), //i
    .p   (dSP_68_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_69 (
    .a   (dSP_69_a[7:0] ), //i
    .d   (dSP_69_d[7:0] ), //i
    .b   (dSP_69_b[7:0] ), //i
    .p   (dSP_69_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_70 (
    .a   (dSP_70_a[7:0] ), //i
    .d   (dSP_70_d[7:0] ), //i
    .b   (dSP_70_b[7:0] ), //i
    .p   (dSP_70_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_71 (
    .a   (dSP_71_a[7:0] ), //i
    .d   (dSP_71_d[7:0] ), //i
    .b   (dSP_71_b[7:0] ), //i
    .p   (dSP_71_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_72 (
    .a   (dSP_72_a[7:0] ), //i
    .d   (dSP_72_d[7:0] ), //i
    .b   (dSP_72_b[7:0] ), //i
    .p   (dSP_72_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_73 (
    .a   (dSP_73_a[7:0] ), //i
    .d   (dSP_73_d[7:0] ), //i
    .b   (dSP_73_b[7:0] ), //i
    .p   (dSP_73_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_74 (
    .a   (dSP_74_a[7:0] ), //i
    .d   (dSP_74_d[7:0] ), //i
    .b   (dSP_74_b[7:0] ), //i
    .p   (dSP_74_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_75 (
    .a   (dSP_75_a[7:0] ), //i
    .d   (dSP_75_d[7:0] ), //i
    .b   (dSP_75_b[7:0] ), //i
    .p   (dSP_75_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_76 (
    .a   (dSP_76_a[7:0] ), //i
    .d   (dSP_76_d[7:0] ), //i
    .b   (dSP_76_b[7:0] ), //i
    .p   (dSP_76_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_77 (
    .a   (dSP_77_a[7:0] ), //i
    .d   (dSP_77_d[7:0] ), //i
    .b   (dSP_77_b[7:0] ), //i
    .p   (dSP_77_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_78 (
    .a   (dSP_78_a[7:0] ), //i
    .d   (dSP_78_d[7:0] ), //i
    .b   (dSP_78_b[7:0] ), //i
    .p   (dSP_78_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_79 (
    .a   (dSP_79_a[7:0] ), //i
    .d   (dSP_79_d[7:0] ), //i
    .b   (dSP_79_b[7:0] ), //i
    .p   (dSP_79_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_80 (
    .a   (dSP_80_a[7:0] ), //i
    .d   (dSP_80_d[7:0] ), //i
    .b   (dSP_80_b[7:0] ), //i
    .p   (dSP_80_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_81 (
    .a   (dSP_81_a[7:0] ), //i
    .d   (dSP_81_d[7:0] ), //i
    .b   (dSP_81_b[7:0] ), //i
    .p   (dSP_81_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_82 (
    .a   (dSP_82_a[7:0] ), //i
    .d   (dSP_82_d[7:0] ), //i
    .b   (dSP_82_b[7:0] ), //i
    .p   (dSP_82_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_83 (
    .a   (dSP_83_a[7:0] ), //i
    .d   (dSP_83_d[7:0] ), //i
    .b   (dSP_83_b[7:0] ), //i
    .p   (dSP_83_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_84 (
    .a   (dSP_84_a[7:0] ), //i
    .d   (dSP_84_d[7:0] ), //i
    .b   (dSP_84_b[7:0] ), //i
    .p   (dSP_84_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_85 (
    .a   (dSP_85_a[7:0] ), //i
    .d   (dSP_85_d[7:0] ), //i
    .b   (dSP_85_b[7:0] ), //i
    .p   (dSP_85_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_86 (
    .a   (dSP_86_a[7:0] ), //i
    .d   (dSP_86_d[7:0] ), //i
    .b   (dSP_86_b[7:0] ), //i
    .p   (dSP_86_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_87 (
    .a   (dSP_87_a[7:0] ), //i
    .d   (dSP_87_d[7:0] ), //i
    .b   (dSP_87_b[7:0] ), //i
    .p   (dSP_87_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_88 (
    .a   (dSP_88_a[7:0] ), //i
    .d   (dSP_88_d[7:0] ), //i
    .b   (dSP_88_b[7:0] ), //i
    .p   (dSP_88_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_89 (
    .a   (dSP_89_a[7:0] ), //i
    .d   (dSP_89_d[7:0] ), //i
    .b   (dSP_89_b[7:0] ), //i
    .p   (dSP_89_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_90 (
    .a   (dSP_90_a[7:0] ), //i
    .d   (dSP_90_d[7:0] ), //i
    .b   (dSP_90_b[7:0] ), //i
    .p   (dSP_90_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_91 (
    .a   (dSP_91_a[7:0] ), //i
    .d   (dSP_91_d[7:0] ), //i
    .b   (dSP_91_b[7:0] ), //i
    .p   (dSP_91_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_92 (
    .a   (dSP_92_a[7:0] ), //i
    .d   (dSP_92_d[7:0] ), //i
    .b   (dSP_92_b[7:0] ), //i
    .p   (dSP_92_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_93 (
    .a   (dSP_93_a[7:0] ), //i
    .d   (dSP_93_d[7:0] ), //i
    .b   (dSP_93_b[7:0] ), //i
    .p   (dSP_93_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_94 (
    .a   (dSP_94_a[7:0] ), //i
    .d   (dSP_94_d[7:0] ), //i
    .b   (dSP_94_b[7:0] ), //i
    .p   (dSP_94_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_95 (
    .a   (dSP_95_a[7:0] ), //i
    .d   (dSP_95_d[7:0] ), //i
    .b   (dSP_95_b[7:0] ), //i
    .p   (dSP_95_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_96 (
    .a   (dSP_96_a[7:0] ), //i
    .d   (dSP_96_d[7:0] ), //i
    .b   (dSP_96_b[7:0] ), //i
    .p   (dSP_96_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_97 (
    .a   (dSP_97_a[7:0] ), //i
    .d   (dSP_97_d[7:0] ), //i
    .b   (dSP_97_b[7:0] ), //i
    .p   (dSP_97_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_98 (
    .a   (dSP_98_a[7:0] ), //i
    .d   (dSP_98_d[7:0] ), //i
    .b   (dSP_98_b[7:0] ), //i
    .p   (dSP_98_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_99 (
    .a   (dSP_99_a[7:0] ), //i
    .d   (dSP_99_d[7:0] ), //i
    .b   (dSP_99_b[7:0] ), //i
    .p   (dSP_99_p[31:0]), //o
    .CLK (clk           )  //i
  );
  DSP dSP_100 (
    .a   (dSP_100_a[7:0] ), //i
    .d   (dSP_100_d[7:0] ), //i
    .b   (dSP_100_b[7:0] ), //i
    .p   (dSP_100_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_101 (
    .a   (dSP_101_a[7:0] ), //i
    .d   (dSP_101_d[7:0] ), //i
    .b   (dSP_101_b[7:0] ), //i
    .p   (dSP_101_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_102 (
    .a   (dSP_102_a[7:0] ), //i
    .d   (dSP_102_d[7:0] ), //i
    .b   (dSP_102_b[7:0] ), //i
    .p   (dSP_102_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_103 (
    .a   (dSP_103_a[7:0] ), //i
    .d   (dSP_103_d[7:0] ), //i
    .b   (dSP_103_b[7:0] ), //i
    .p   (dSP_103_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_104 (
    .a   (dSP_104_a[7:0] ), //i
    .d   (dSP_104_d[7:0] ), //i
    .b   (dSP_104_b[7:0] ), //i
    .p   (dSP_104_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_105 (
    .a   (dSP_105_a[7:0] ), //i
    .d   (dSP_105_d[7:0] ), //i
    .b   (dSP_105_b[7:0] ), //i
    .p   (dSP_105_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_106 (
    .a   (dSP_106_a[7:0] ), //i
    .d   (dSP_106_d[7:0] ), //i
    .b   (dSP_106_b[7:0] ), //i
    .p   (dSP_106_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_107 (
    .a   (dSP_107_a[7:0] ), //i
    .d   (dSP_107_d[7:0] ), //i
    .b   (dSP_107_b[7:0] ), //i
    .p   (dSP_107_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_108 (
    .a   (dSP_108_a[7:0] ), //i
    .d   (dSP_108_d[7:0] ), //i
    .b   (dSP_108_b[7:0] ), //i
    .p   (dSP_108_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_109 (
    .a   (dSP_109_a[7:0] ), //i
    .d   (dSP_109_d[7:0] ), //i
    .b   (dSP_109_b[7:0] ), //i
    .p   (dSP_109_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_110 (
    .a   (dSP_110_a[7:0] ), //i
    .d   (dSP_110_d[7:0] ), //i
    .b   (dSP_110_b[7:0] ), //i
    .p   (dSP_110_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_111 (
    .a   (dSP_111_a[7:0] ), //i
    .d   (dSP_111_d[7:0] ), //i
    .b   (dSP_111_b[7:0] ), //i
    .p   (dSP_111_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_112 (
    .a   (dSP_112_a[7:0] ), //i
    .d   (dSP_112_d[7:0] ), //i
    .b   (dSP_112_b[7:0] ), //i
    .p   (dSP_112_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_113 (
    .a   (dSP_113_a[7:0] ), //i
    .d   (dSP_113_d[7:0] ), //i
    .b   (dSP_113_b[7:0] ), //i
    .p   (dSP_113_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_114 (
    .a   (dSP_114_a[7:0] ), //i
    .d   (dSP_114_d[7:0] ), //i
    .b   (dSP_114_b[7:0] ), //i
    .p   (dSP_114_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_115 (
    .a   (dSP_115_a[7:0] ), //i
    .d   (dSP_115_d[7:0] ), //i
    .b   (dSP_115_b[7:0] ), //i
    .p   (dSP_115_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_116 (
    .a   (dSP_116_a[7:0] ), //i
    .d   (dSP_116_d[7:0] ), //i
    .b   (dSP_116_b[7:0] ), //i
    .p   (dSP_116_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_117 (
    .a   (dSP_117_a[7:0] ), //i
    .d   (dSP_117_d[7:0] ), //i
    .b   (dSP_117_b[7:0] ), //i
    .p   (dSP_117_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_118 (
    .a   (dSP_118_a[7:0] ), //i
    .d   (dSP_118_d[7:0] ), //i
    .b   (dSP_118_b[7:0] ), //i
    .p   (dSP_118_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_119 (
    .a   (dSP_119_a[7:0] ), //i
    .d   (dSP_119_d[7:0] ), //i
    .b   (dSP_119_b[7:0] ), //i
    .p   (dSP_119_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_120 (
    .a   (dSP_120_a[7:0] ), //i
    .d   (dSP_120_d[7:0] ), //i
    .b   (dSP_120_b[7:0] ), //i
    .p   (dSP_120_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_121 (
    .a   (dSP_121_a[7:0] ), //i
    .d   (dSP_121_d[7:0] ), //i
    .b   (dSP_121_b[7:0] ), //i
    .p   (dSP_121_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_122 (
    .a   (dSP_122_a[7:0] ), //i
    .d   (dSP_122_d[7:0] ), //i
    .b   (dSP_122_b[7:0] ), //i
    .p   (dSP_122_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_123 (
    .a   (dSP_123_a[7:0] ), //i
    .d   (dSP_123_d[7:0] ), //i
    .b   (dSP_123_b[7:0] ), //i
    .p   (dSP_123_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_124 (
    .a   (dSP_124_a[7:0] ), //i
    .d   (dSP_124_d[7:0] ), //i
    .b   (dSP_124_b[7:0] ), //i
    .p   (dSP_124_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_125 (
    .a   (dSP_125_a[7:0] ), //i
    .d   (dSP_125_d[7:0] ), //i
    .b   (dSP_125_b[7:0] ), //i
    .p   (dSP_125_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_126 (
    .a   (dSP_126_a[7:0] ), //i
    .d   (dSP_126_d[7:0] ), //i
    .b   (dSP_126_b[7:0] ), //i
    .p   (dSP_126_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_127 (
    .a   (dSP_127_a[7:0] ), //i
    .d   (dSP_127_d[7:0] ), //i
    .b   (dSP_127_b[7:0] ), //i
    .p   (dSP_127_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_128 (
    .a   (dSP_128_a[7:0] ), //i
    .d   (dSP_128_d[7:0] ), //i
    .b   (dSP_128_b[7:0] ), //i
    .p   (dSP_128_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_129 (
    .a   (dSP_129_a[7:0] ), //i
    .d   (dSP_129_d[7:0] ), //i
    .b   (dSP_129_b[7:0] ), //i
    .p   (dSP_129_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_130 (
    .a   (dSP_130_a[7:0] ), //i
    .d   (dSP_130_d[7:0] ), //i
    .b   (dSP_130_b[7:0] ), //i
    .p   (dSP_130_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_131 (
    .a   (dSP_131_a[7:0] ), //i
    .d   (dSP_131_d[7:0] ), //i
    .b   (dSP_131_b[7:0] ), //i
    .p   (dSP_131_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_132 (
    .a   (dSP_132_a[7:0] ), //i
    .d   (dSP_132_d[7:0] ), //i
    .b   (dSP_132_b[7:0] ), //i
    .p   (dSP_132_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_133 (
    .a   (dSP_133_a[7:0] ), //i
    .d   (dSP_133_d[7:0] ), //i
    .b   (dSP_133_b[7:0] ), //i
    .p   (dSP_133_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_134 (
    .a   (dSP_134_a[7:0] ), //i
    .d   (dSP_134_d[7:0] ), //i
    .b   (dSP_134_b[7:0] ), //i
    .p   (dSP_134_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_135 (
    .a   (dSP_135_a[7:0] ), //i
    .d   (dSP_135_d[7:0] ), //i
    .b   (dSP_135_b[7:0] ), //i
    .p   (dSP_135_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_136 (
    .a   (dSP_136_a[7:0] ), //i
    .d   (dSP_136_d[7:0] ), //i
    .b   (dSP_136_b[7:0] ), //i
    .p   (dSP_136_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_137 (
    .a   (dSP_137_a[7:0] ), //i
    .d   (dSP_137_d[7:0] ), //i
    .b   (dSP_137_b[7:0] ), //i
    .p   (dSP_137_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_138 (
    .a   (dSP_138_a[7:0] ), //i
    .d   (dSP_138_d[7:0] ), //i
    .b   (dSP_138_b[7:0] ), //i
    .p   (dSP_138_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_139 (
    .a   (dSP_139_a[7:0] ), //i
    .d   (dSP_139_d[7:0] ), //i
    .b   (dSP_139_b[7:0] ), //i
    .p   (dSP_139_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_140 (
    .a   (dSP_140_a[7:0] ), //i
    .d   (dSP_140_d[7:0] ), //i
    .b   (dSP_140_b[7:0] ), //i
    .p   (dSP_140_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_141 (
    .a   (dSP_141_a[7:0] ), //i
    .d   (dSP_141_d[7:0] ), //i
    .b   (dSP_141_b[7:0] ), //i
    .p   (dSP_141_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_142 (
    .a   (dSP_142_a[7:0] ), //i
    .d   (dSP_142_d[7:0] ), //i
    .b   (dSP_142_b[7:0] ), //i
    .p   (dSP_142_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_143 (
    .a   (dSP_143_a[7:0] ), //i
    .d   (dSP_143_d[7:0] ), //i
    .b   (dSP_143_b[7:0] ), //i
    .p   (dSP_143_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_144 (
    .a   (dSP_144_a[7:0] ), //i
    .d   (dSP_144_d[7:0] ), //i
    .b   (dSP_144_b[7:0] ), //i
    .p   (dSP_144_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_145 (
    .a   (dSP_145_a[7:0] ), //i
    .d   (dSP_145_d[7:0] ), //i
    .b   (dSP_145_b[7:0] ), //i
    .p   (dSP_145_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_146 (
    .a   (dSP_146_a[7:0] ), //i
    .d   (dSP_146_d[7:0] ), //i
    .b   (dSP_146_b[7:0] ), //i
    .p   (dSP_146_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_147 (
    .a   (dSP_147_a[7:0] ), //i
    .d   (dSP_147_d[7:0] ), //i
    .b   (dSP_147_b[7:0] ), //i
    .p   (dSP_147_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_148 (
    .a   (dSP_148_a[7:0] ), //i
    .d   (dSP_148_d[7:0] ), //i
    .b   (dSP_148_b[7:0] ), //i
    .p   (dSP_148_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_149 (
    .a   (dSP_149_a[7:0] ), //i
    .d   (dSP_149_d[7:0] ), //i
    .b   (dSP_149_b[7:0] ), //i
    .p   (dSP_149_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_150 (
    .a   (dSP_150_a[7:0] ), //i
    .d   (dSP_150_d[7:0] ), //i
    .b   (dSP_150_b[7:0] ), //i
    .p   (dSP_150_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_151 (
    .a   (dSP_151_a[7:0] ), //i
    .d   (dSP_151_d[7:0] ), //i
    .b   (dSP_151_b[7:0] ), //i
    .p   (dSP_151_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_152 (
    .a   (dSP_152_a[7:0] ), //i
    .d   (dSP_152_d[7:0] ), //i
    .b   (dSP_152_b[7:0] ), //i
    .p   (dSP_152_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_153 (
    .a   (dSP_153_a[7:0] ), //i
    .d   (dSP_153_d[7:0] ), //i
    .b   (dSP_153_b[7:0] ), //i
    .p   (dSP_153_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_154 (
    .a   (dSP_154_a[7:0] ), //i
    .d   (dSP_154_d[7:0] ), //i
    .b   (dSP_154_b[7:0] ), //i
    .p   (dSP_154_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_155 (
    .a   (dSP_155_a[7:0] ), //i
    .d   (dSP_155_d[7:0] ), //i
    .b   (dSP_155_b[7:0] ), //i
    .p   (dSP_155_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_156 (
    .a   (dSP_156_a[7:0] ), //i
    .d   (dSP_156_d[7:0] ), //i
    .b   (dSP_156_b[7:0] ), //i
    .p   (dSP_156_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_157 (
    .a   (dSP_157_a[7:0] ), //i
    .d   (dSP_157_d[7:0] ), //i
    .b   (dSP_157_b[7:0] ), //i
    .p   (dSP_157_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_158 (
    .a   (dSP_158_a[7:0] ), //i
    .d   (dSP_158_d[7:0] ), //i
    .b   (dSP_158_b[7:0] ), //i
    .p   (dSP_158_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_159 (
    .a   (dSP_159_a[7:0] ), //i
    .d   (dSP_159_d[7:0] ), //i
    .b   (dSP_159_b[7:0] ), //i
    .p   (dSP_159_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_160 (
    .a   (dSP_160_a[7:0] ), //i
    .d   (dSP_160_d[7:0] ), //i
    .b   (dSP_160_b[7:0] ), //i
    .p   (dSP_160_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_161 (
    .a   (dSP_161_a[7:0] ), //i
    .d   (dSP_161_d[7:0] ), //i
    .b   (dSP_161_b[7:0] ), //i
    .p   (dSP_161_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_162 (
    .a   (dSP_162_a[7:0] ), //i
    .d   (dSP_162_d[7:0] ), //i
    .b   (dSP_162_b[7:0] ), //i
    .p   (dSP_162_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_163 (
    .a   (dSP_163_a[7:0] ), //i
    .d   (dSP_163_d[7:0] ), //i
    .b   (dSP_163_b[7:0] ), //i
    .p   (dSP_163_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_164 (
    .a   (dSP_164_a[7:0] ), //i
    .d   (dSP_164_d[7:0] ), //i
    .b   (dSP_164_b[7:0] ), //i
    .p   (dSP_164_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_165 (
    .a   (dSP_165_a[7:0] ), //i
    .d   (dSP_165_d[7:0] ), //i
    .b   (dSP_165_b[7:0] ), //i
    .p   (dSP_165_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_166 (
    .a   (dSP_166_a[7:0] ), //i
    .d   (dSP_166_d[7:0] ), //i
    .b   (dSP_166_b[7:0] ), //i
    .p   (dSP_166_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_167 (
    .a   (dSP_167_a[7:0] ), //i
    .d   (dSP_167_d[7:0] ), //i
    .b   (dSP_167_b[7:0] ), //i
    .p   (dSP_167_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_168 (
    .a   (dSP_168_a[7:0] ), //i
    .d   (dSP_168_d[7:0] ), //i
    .b   (dSP_168_b[7:0] ), //i
    .p   (dSP_168_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_169 (
    .a   (dSP_169_a[7:0] ), //i
    .d   (dSP_169_d[7:0] ), //i
    .b   (dSP_169_b[7:0] ), //i
    .p   (dSP_169_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_170 (
    .a   (dSP_170_a[7:0] ), //i
    .d   (dSP_170_d[7:0] ), //i
    .b   (dSP_170_b[7:0] ), //i
    .p   (dSP_170_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_171 (
    .a   (dSP_171_a[7:0] ), //i
    .d   (dSP_171_d[7:0] ), //i
    .b   (dSP_171_b[7:0] ), //i
    .p   (dSP_171_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_172 (
    .a   (dSP_172_a[7:0] ), //i
    .d   (dSP_172_d[7:0] ), //i
    .b   (dSP_172_b[7:0] ), //i
    .p   (dSP_172_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_173 (
    .a   (dSP_173_a[7:0] ), //i
    .d   (dSP_173_d[7:0] ), //i
    .b   (dSP_173_b[7:0] ), //i
    .p   (dSP_173_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_174 (
    .a   (dSP_174_a[7:0] ), //i
    .d   (dSP_174_d[7:0] ), //i
    .b   (dSP_174_b[7:0] ), //i
    .p   (dSP_174_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_175 (
    .a   (dSP_175_a[7:0] ), //i
    .d   (dSP_175_d[7:0] ), //i
    .b   (dSP_175_b[7:0] ), //i
    .p   (dSP_175_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_176 (
    .a   (dSP_176_a[7:0] ), //i
    .d   (dSP_176_d[7:0] ), //i
    .b   (dSP_176_b[7:0] ), //i
    .p   (dSP_176_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_177 (
    .a   (dSP_177_a[7:0] ), //i
    .d   (dSP_177_d[7:0] ), //i
    .b   (dSP_177_b[7:0] ), //i
    .p   (dSP_177_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_178 (
    .a   (dSP_178_a[7:0] ), //i
    .d   (dSP_178_d[7:0] ), //i
    .b   (dSP_178_b[7:0] ), //i
    .p   (dSP_178_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_179 (
    .a   (dSP_179_a[7:0] ), //i
    .d   (dSP_179_d[7:0] ), //i
    .b   (dSP_179_b[7:0] ), //i
    .p   (dSP_179_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_180 (
    .a   (dSP_180_a[7:0] ), //i
    .d   (dSP_180_d[7:0] ), //i
    .b   (dSP_180_b[7:0] ), //i
    .p   (dSP_180_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_181 (
    .a   (dSP_181_a[7:0] ), //i
    .d   (dSP_181_d[7:0] ), //i
    .b   (dSP_181_b[7:0] ), //i
    .p   (dSP_181_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_182 (
    .a   (dSP_182_a[7:0] ), //i
    .d   (dSP_182_d[7:0] ), //i
    .b   (dSP_182_b[7:0] ), //i
    .p   (dSP_182_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_183 (
    .a   (dSP_183_a[7:0] ), //i
    .d   (dSP_183_d[7:0] ), //i
    .b   (dSP_183_b[7:0] ), //i
    .p   (dSP_183_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_184 (
    .a   (dSP_184_a[7:0] ), //i
    .d   (dSP_184_d[7:0] ), //i
    .b   (dSP_184_b[7:0] ), //i
    .p   (dSP_184_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_185 (
    .a   (dSP_185_a[7:0] ), //i
    .d   (dSP_185_d[7:0] ), //i
    .b   (dSP_185_b[7:0] ), //i
    .p   (dSP_185_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_186 (
    .a   (dSP_186_a[7:0] ), //i
    .d   (dSP_186_d[7:0] ), //i
    .b   (dSP_186_b[7:0] ), //i
    .p   (dSP_186_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_187 (
    .a   (dSP_187_a[7:0] ), //i
    .d   (dSP_187_d[7:0] ), //i
    .b   (dSP_187_b[7:0] ), //i
    .p   (dSP_187_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_188 (
    .a   (dSP_188_a[7:0] ), //i
    .d   (dSP_188_d[7:0] ), //i
    .b   (dSP_188_b[7:0] ), //i
    .p   (dSP_188_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_189 (
    .a   (dSP_189_a[7:0] ), //i
    .d   (dSP_189_d[7:0] ), //i
    .b   (dSP_189_b[7:0] ), //i
    .p   (dSP_189_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_190 (
    .a   (dSP_190_a[7:0] ), //i
    .d   (dSP_190_d[7:0] ), //i
    .b   (dSP_190_b[7:0] ), //i
    .p   (dSP_190_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_191 (
    .a   (dSP_191_a[7:0] ), //i
    .d   (dSP_191_d[7:0] ), //i
    .b   (dSP_191_b[7:0] ), //i
    .p   (dSP_191_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_192 (
    .a   (dSP_192_a[7:0] ), //i
    .d   (dSP_192_d[7:0] ), //i
    .b   (dSP_192_b[7:0] ), //i
    .p   (dSP_192_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_193 (
    .a   (dSP_193_a[7:0] ), //i
    .d   (dSP_193_d[7:0] ), //i
    .b   (dSP_193_b[7:0] ), //i
    .p   (dSP_193_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_194 (
    .a   (dSP_194_a[7:0] ), //i
    .d   (dSP_194_d[7:0] ), //i
    .b   (dSP_194_b[7:0] ), //i
    .p   (dSP_194_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_195 (
    .a   (dSP_195_a[7:0] ), //i
    .d   (dSP_195_d[7:0] ), //i
    .b   (dSP_195_b[7:0] ), //i
    .p   (dSP_195_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_196 (
    .a   (dSP_196_a[7:0] ), //i
    .d   (dSP_196_d[7:0] ), //i
    .b   (dSP_196_b[7:0] ), //i
    .p   (dSP_196_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_197 (
    .a   (dSP_197_a[7:0] ), //i
    .d   (dSP_197_d[7:0] ), //i
    .b   (dSP_197_b[7:0] ), //i
    .p   (dSP_197_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_198 (
    .a   (dSP_198_a[7:0] ), //i
    .d   (dSP_198_d[7:0] ), //i
    .b   (dSP_198_b[7:0] ), //i
    .p   (dSP_198_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_199 (
    .a   (dSP_199_a[7:0] ), //i
    .d   (dSP_199_d[7:0] ), //i
    .b   (dSP_199_b[7:0] ), //i
    .p   (dSP_199_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_200 (
    .a   (dSP_200_a[7:0] ), //i
    .d   (dSP_200_d[7:0] ), //i
    .b   (dSP_200_b[7:0] ), //i
    .p   (dSP_200_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_201 (
    .a   (dSP_201_a[7:0] ), //i
    .d   (dSP_201_d[7:0] ), //i
    .b   (dSP_201_b[7:0] ), //i
    .p   (dSP_201_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_202 (
    .a   (dSP_202_a[7:0] ), //i
    .d   (dSP_202_d[7:0] ), //i
    .b   (dSP_202_b[7:0] ), //i
    .p   (dSP_202_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_203 (
    .a   (dSP_203_a[7:0] ), //i
    .d   (dSP_203_d[7:0] ), //i
    .b   (dSP_203_b[7:0] ), //i
    .p   (dSP_203_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_204 (
    .a   (dSP_204_a[7:0] ), //i
    .d   (dSP_204_d[7:0] ), //i
    .b   (dSP_204_b[7:0] ), //i
    .p   (dSP_204_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_205 (
    .a   (dSP_205_a[7:0] ), //i
    .d   (dSP_205_d[7:0] ), //i
    .b   (dSP_205_b[7:0] ), //i
    .p   (dSP_205_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_206 (
    .a   (dSP_206_a[7:0] ), //i
    .d   (dSP_206_d[7:0] ), //i
    .b   (dSP_206_b[7:0] ), //i
    .p   (dSP_206_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_207 (
    .a   (dSP_207_a[7:0] ), //i
    .d   (dSP_207_d[7:0] ), //i
    .b   (dSP_207_b[7:0] ), //i
    .p   (dSP_207_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_208 (
    .a   (dSP_208_a[7:0] ), //i
    .d   (dSP_208_d[7:0] ), //i
    .b   (dSP_208_b[7:0] ), //i
    .p   (dSP_208_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_209 (
    .a   (dSP_209_a[7:0] ), //i
    .d   (dSP_209_d[7:0] ), //i
    .b   (dSP_209_b[7:0] ), //i
    .p   (dSP_209_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_210 (
    .a   (dSP_210_a[7:0] ), //i
    .d   (dSP_210_d[7:0] ), //i
    .b   (dSP_210_b[7:0] ), //i
    .p   (dSP_210_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_211 (
    .a   (dSP_211_a[7:0] ), //i
    .d   (dSP_211_d[7:0] ), //i
    .b   (dSP_211_b[7:0] ), //i
    .p   (dSP_211_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_212 (
    .a   (dSP_212_a[7:0] ), //i
    .d   (dSP_212_d[7:0] ), //i
    .b   (dSP_212_b[7:0] ), //i
    .p   (dSP_212_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_213 (
    .a   (dSP_213_a[7:0] ), //i
    .d   (dSP_213_d[7:0] ), //i
    .b   (dSP_213_b[7:0] ), //i
    .p   (dSP_213_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_214 (
    .a   (dSP_214_a[7:0] ), //i
    .d   (dSP_214_d[7:0] ), //i
    .b   (dSP_214_b[7:0] ), //i
    .p   (dSP_214_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_215 (
    .a   (dSP_215_a[7:0] ), //i
    .d   (dSP_215_d[7:0] ), //i
    .b   (dSP_215_b[7:0] ), //i
    .p   (dSP_215_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_216 (
    .a   (dSP_216_a[7:0] ), //i
    .d   (dSP_216_d[7:0] ), //i
    .b   (dSP_216_b[7:0] ), //i
    .p   (dSP_216_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_217 (
    .a   (dSP_217_a[7:0] ), //i
    .d   (dSP_217_d[7:0] ), //i
    .b   (dSP_217_b[7:0] ), //i
    .p   (dSP_217_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_218 (
    .a   (dSP_218_a[7:0] ), //i
    .d   (dSP_218_d[7:0] ), //i
    .b   (dSP_218_b[7:0] ), //i
    .p   (dSP_218_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_219 (
    .a   (dSP_219_a[7:0] ), //i
    .d   (dSP_219_d[7:0] ), //i
    .b   (dSP_219_b[7:0] ), //i
    .p   (dSP_219_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_220 (
    .a   (dSP_220_a[7:0] ), //i
    .d   (dSP_220_d[7:0] ), //i
    .b   (dSP_220_b[7:0] ), //i
    .p   (dSP_220_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_221 (
    .a   (dSP_221_a[7:0] ), //i
    .d   (dSP_221_d[7:0] ), //i
    .b   (dSP_221_b[7:0] ), //i
    .p   (dSP_221_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_222 (
    .a   (dSP_222_a[7:0] ), //i
    .d   (dSP_222_d[7:0] ), //i
    .b   (dSP_222_b[7:0] ), //i
    .p   (dSP_222_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_223 (
    .a   (dSP_223_a[7:0] ), //i
    .d   (dSP_223_d[7:0] ), //i
    .b   (dSP_223_b[7:0] ), //i
    .p   (dSP_223_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_224 (
    .a   (dSP_224_a[7:0] ), //i
    .d   (dSP_224_d[7:0] ), //i
    .b   (dSP_224_b[7:0] ), //i
    .p   (dSP_224_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_225 (
    .a   (dSP_225_a[7:0] ), //i
    .d   (dSP_225_d[7:0] ), //i
    .b   (dSP_225_b[7:0] ), //i
    .p   (dSP_225_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_226 (
    .a   (dSP_226_a[7:0] ), //i
    .d   (dSP_226_d[7:0] ), //i
    .b   (dSP_226_b[7:0] ), //i
    .p   (dSP_226_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_227 (
    .a   (dSP_227_a[7:0] ), //i
    .d   (dSP_227_d[7:0] ), //i
    .b   (dSP_227_b[7:0] ), //i
    .p   (dSP_227_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_228 (
    .a   (dSP_228_a[7:0] ), //i
    .d   (dSP_228_d[7:0] ), //i
    .b   (dSP_228_b[7:0] ), //i
    .p   (dSP_228_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_229 (
    .a   (dSP_229_a[7:0] ), //i
    .d   (dSP_229_d[7:0] ), //i
    .b   (dSP_229_b[7:0] ), //i
    .p   (dSP_229_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_230 (
    .a   (dSP_230_a[7:0] ), //i
    .d   (dSP_230_d[7:0] ), //i
    .b   (dSP_230_b[7:0] ), //i
    .p   (dSP_230_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_231 (
    .a   (dSP_231_a[7:0] ), //i
    .d   (dSP_231_d[7:0] ), //i
    .b   (dSP_231_b[7:0] ), //i
    .p   (dSP_231_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_232 (
    .a   (dSP_232_a[7:0] ), //i
    .d   (dSP_232_d[7:0] ), //i
    .b   (dSP_232_b[7:0] ), //i
    .p   (dSP_232_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_233 (
    .a   (dSP_233_a[7:0] ), //i
    .d   (dSP_233_d[7:0] ), //i
    .b   (dSP_233_b[7:0] ), //i
    .p   (dSP_233_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_234 (
    .a   (dSP_234_a[7:0] ), //i
    .d   (dSP_234_d[7:0] ), //i
    .b   (dSP_234_b[7:0] ), //i
    .p   (dSP_234_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_235 (
    .a   (dSP_235_a[7:0] ), //i
    .d   (dSP_235_d[7:0] ), //i
    .b   (dSP_235_b[7:0] ), //i
    .p   (dSP_235_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_236 (
    .a   (dSP_236_a[7:0] ), //i
    .d   (dSP_236_d[7:0] ), //i
    .b   (dSP_236_b[7:0] ), //i
    .p   (dSP_236_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_237 (
    .a   (dSP_237_a[7:0] ), //i
    .d   (dSP_237_d[7:0] ), //i
    .b   (dSP_237_b[7:0] ), //i
    .p   (dSP_237_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_238 (
    .a   (dSP_238_a[7:0] ), //i
    .d   (dSP_238_d[7:0] ), //i
    .b   (dSP_238_b[7:0] ), //i
    .p   (dSP_238_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_239 (
    .a   (dSP_239_a[7:0] ), //i
    .d   (dSP_239_d[7:0] ), //i
    .b   (dSP_239_b[7:0] ), //i
    .p   (dSP_239_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_240 (
    .a   (dSP_240_a[7:0] ), //i
    .d   (dSP_240_d[7:0] ), //i
    .b   (dSP_240_b[7:0] ), //i
    .p   (dSP_240_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_241 (
    .a   (dSP_241_a[7:0] ), //i
    .d   (dSP_241_d[7:0] ), //i
    .b   (dSP_241_b[7:0] ), //i
    .p   (dSP_241_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_242 (
    .a   (dSP_242_a[7:0] ), //i
    .d   (dSP_242_d[7:0] ), //i
    .b   (dSP_242_b[7:0] ), //i
    .p   (dSP_242_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_243 (
    .a   (dSP_243_a[7:0] ), //i
    .d   (dSP_243_d[7:0] ), //i
    .b   (dSP_243_b[7:0] ), //i
    .p   (dSP_243_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_244 (
    .a   (dSP_244_a[7:0] ), //i
    .d   (dSP_244_d[7:0] ), //i
    .b   (dSP_244_b[7:0] ), //i
    .p   (dSP_244_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_245 (
    .a   (dSP_245_a[7:0] ), //i
    .d   (dSP_245_d[7:0] ), //i
    .b   (dSP_245_b[7:0] ), //i
    .p   (dSP_245_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_246 (
    .a   (dSP_246_a[7:0] ), //i
    .d   (dSP_246_d[7:0] ), //i
    .b   (dSP_246_b[7:0] ), //i
    .p   (dSP_246_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_247 (
    .a   (dSP_247_a[7:0] ), //i
    .d   (dSP_247_d[7:0] ), //i
    .b   (dSP_247_b[7:0] ), //i
    .p   (dSP_247_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_248 (
    .a   (dSP_248_a[7:0] ), //i
    .d   (dSP_248_d[7:0] ), //i
    .b   (dSP_248_b[7:0] ), //i
    .p   (dSP_248_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_249 (
    .a   (dSP_249_a[7:0] ), //i
    .d   (dSP_249_d[7:0] ), //i
    .b   (dSP_249_b[7:0] ), //i
    .p   (dSP_249_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_250 (
    .a   (dSP_250_a[7:0] ), //i
    .d   (dSP_250_d[7:0] ), //i
    .b   (dSP_250_b[7:0] ), //i
    .p   (dSP_250_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_251 (
    .a   (dSP_251_a[7:0] ), //i
    .d   (dSP_251_d[7:0] ), //i
    .b   (dSP_251_b[7:0] ), //i
    .p   (dSP_251_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_252 (
    .a   (dSP_252_a[7:0] ), //i
    .d   (dSP_252_d[7:0] ), //i
    .b   (dSP_252_b[7:0] ), //i
    .p   (dSP_252_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_253 (
    .a   (dSP_253_a[7:0] ), //i
    .d   (dSP_253_d[7:0] ), //i
    .b   (dSP_253_b[7:0] ), //i
    .p   (dSP_253_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_254 (
    .a   (dSP_254_a[7:0] ), //i
    .d   (dSP_254_d[7:0] ), //i
    .b   (dSP_254_b[7:0] ), //i
    .p   (dSP_254_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_255 (
    .a   (dSP_255_a[7:0] ), //i
    .d   (dSP_255_d[7:0] ), //i
    .b   (dSP_255_b[7:0] ), //i
    .p   (dSP_255_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_256 (
    .a   (dSP_256_a[7:0] ), //i
    .d   (dSP_256_d[7:0] ), //i
    .b   (dSP_256_b[7:0] ), //i
    .p   (dSP_256_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_257 (
    .a   (dSP_257_a[7:0] ), //i
    .d   (dSP_257_d[7:0] ), //i
    .b   (dSP_257_b[7:0] ), //i
    .p   (dSP_257_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_258 (
    .a   (dSP_258_a[7:0] ), //i
    .d   (dSP_258_d[7:0] ), //i
    .b   (dSP_258_b[7:0] ), //i
    .p   (dSP_258_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_259 (
    .a   (dSP_259_a[7:0] ), //i
    .d   (dSP_259_d[7:0] ), //i
    .b   (dSP_259_b[7:0] ), //i
    .p   (dSP_259_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_260 (
    .a   (dSP_260_a[7:0] ), //i
    .d   (dSP_260_d[7:0] ), //i
    .b   (dSP_260_b[7:0] ), //i
    .p   (dSP_260_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_261 (
    .a   (dSP_261_a[7:0] ), //i
    .d   (dSP_261_d[7:0] ), //i
    .b   (dSP_261_b[7:0] ), //i
    .p   (dSP_261_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_262 (
    .a   (dSP_262_a[7:0] ), //i
    .d   (dSP_262_d[7:0] ), //i
    .b   (dSP_262_b[7:0] ), //i
    .p   (dSP_262_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_263 (
    .a   (dSP_263_a[7:0] ), //i
    .d   (dSP_263_d[7:0] ), //i
    .b   (dSP_263_b[7:0] ), //i
    .p   (dSP_263_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_264 (
    .a   (dSP_264_a[7:0] ), //i
    .d   (dSP_264_d[7:0] ), //i
    .b   (dSP_264_b[7:0] ), //i
    .p   (dSP_264_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_265 (
    .a   (dSP_265_a[7:0] ), //i
    .d   (dSP_265_d[7:0] ), //i
    .b   (dSP_265_b[7:0] ), //i
    .p   (dSP_265_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_266 (
    .a   (dSP_266_a[7:0] ), //i
    .d   (dSP_266_d[7:0] ), //i
    .b   (dSP_266_b[7:0] ), //i
    .p   (dSP_266_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_267 (
    .a   (dSP_267_a[7:0] ), //i
    .d   (dSP_267_d[7:0] ), //i
    .b   (dSP_267_b[7:0] ), //i
    .p   (dSP_267_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_268 (
    .a   (dSP_268_a[7:0] ), //i
    .d   (dSP_268_d[7:0] ), //i
    .b   (dSP_268_b[7:0] ), //i
    .p   (dSP_268_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_269 (
    .a   (dSP_269_a[7:0] ), //i
    .d   (dSP_269_d[7:0] ), //i
    .b   (dSP_269_b[7:0] ), //i
    .p   (dSP_269_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_270 (
    .a   (dSP_270_a[7:0] ), //i
    .d   (dSP_270_d[7:0] ), //i
    .b   (dSP_270_b[7:0] ), //i
    .p   (dSP_270_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_271 (
    .a   (dSP_271_a[7:0] ), //i
    .d   (dSP_271_d[7:0] ), //i
    .b   (dSP_271_b[7:0] ), //i
    .p   (dSP_271_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_272 (
    .a   (dSP_272_a[7:0] ), //i
    .d   (dSP_272_d[7:0] ), //i
    .b   (dSP_272_b[7:0] ), //i
    .p   (dSP_272_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_273 (
    .a   (dSP_273_a[7:0] ), //i
    .d   (dSP_273_d[7:0] ), //i
    .b   (dSP_273_b[7:0] ), //i
    .p   (dSP_273_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_274 (
    .a   (dSP_274_a[7:0] ), //i
    .d   (dSP_274_d[7:0] ), //i
    .b   (dSP_274_b[7:0] ), //i
    .p   (dSP_274_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_275 (
    .a   (dSP_275_a[7:0] ), //i
    .d   (dSP_275_d[7:0] ), //i
    .b   (dSP_275_b[7:0] ), //i
    .p   (dSP_275_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_276 (
    .a   (dSP_276_a[7:0] ), //i
    .d   (dSP_276_d[7:0] ), //i
    .b   (dSP_276_b[7:0] ), //i
    .p   (dSP_276_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_277 (
    .a   (dSP_277_a[7:0] ), //i
    .d   (dSP_277_d[7:0] ), //i
    .b   (dSP_277_b[7:0] ), //i
    .p   (dSP_277_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_278 (
    .a   (dSP_278_a[7:0] ), //i
    .d   (dSP_278_d[7:0] ), //i
    .b   (dSP_278_b[7:0] ), //i
    .p   (dSP_278_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_279 (
    .a   (dSP_279_a[7:0] ), //i
    .d   (dSP_279_d[7:0] ), //i
    .b   (dSP_279_b[7:0] ), //i
    .p   (dSP_279_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_280 (
    .a   (dSP_280_a[7:0] ), //i
    .d   (dSP_280_d[7:0] ), //i
    .b   (dSP_280_b[7:0] ), //i
    .p   (dSP_280_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_281 (
    .a   (dSP_281_a[7:0] ), //i
    .d   (dSP_281_d[7:0] ), //i
    .b   (dSP_281_b[7:0] ), //i
    .p   (dSP_281_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_282 (
    .a   (dSP_282_a[7:0] ), //i
    .d   (dSP_282_d[7:0] ), //i
    .b   (dSP_282_b[7:0] ), //i
    .p   (dSP_282_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_283 (
    .a   (dSP_283_a[7:0] ), //i
    .d   (dSP_283_d[7:0] ), //i
    .b   (dSP_283_b[7:0] ), //i
    .p   (dSP_283_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_284 (
    .a   (dSP_284_a[7:0] ), //i
    .d   (dSP_284_d[7:0] ), //i
    .b   (dSP_284_b[7:0] ), //i
    .p   (dSP_284_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_285 (
    .a   (dSP_285_a[7:0] ), //i
    .d   (dSP_285_d[7:0] ), //i
    .b   (dSP_285_b[7:0] ), //i
    .p   (dSP_285_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_286 (
    .a   (dSP_286_a[7:0] ), //i
    .d   (dSP_286_d[7:0] ), //i
    .b   (dSP_286_b[7:0] ), //i
    .p   (dSP_286_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_287 (
    .a   (dSP_287_a[7:0] ), //i
    .d   (dSP_287_d[7:0] ), //i
    .b   (dSP_287_b[7:0] ), //i
    .p   (dSP_287_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_288 (
    .a   (dSP_288_a[7:0] ), //i
    .d   (dSP_288_d[7:0] ), //i
    .b   (dSP_288_b[7:0] ), //i
    .p   (dSP_288_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_289 (
    .a   (dSP_289_a[7:0] ), //i
    .d   (dSP_289_d[7:0] ), //i
    .b   (dSP_289_b[7:0] ), //i
    .p   (dSP_289_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_290 (
    .a   (dSP_290_a[7:0] ), //i
    .d   (dSP_290_d[7:0] ), //i
    .b   (dSP_290_b[7:0] ), //i
    .p   (dSP_290_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_291 (
    .a   (dSP_291_a[7:0] ), //i
    .d   (dSP_291_d[7:0] ), //i
    .b   (dSP_291_b[7:0] ), //i
    .p   (dSP_291_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_292 (
    .a   (dSP_292_a[7:0] ), //i
    .d   (dSP_292_d[7:0] ), //i
    .b   (dSP_292_b[7:0] ), //i
    .p   (dSP_292_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_293 (
    .a   (dSP_293_a[7:0] ), //i
    .d   (dSP_293_d[7:0] ), //i
    .b   (dSP_293_b[7:0] ), //i
    .p   (dSP_293_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_294 (
    .a   (dSP_294_a[7:0] ), //i
    .d   (dSP_294_d[7:0] ), //i
    .b   (dSP_294_b[7:0] ), //i
    .p   (dSP_294_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_295 (
    .a   (dSP_295_a[7:0] ), //i
    .d   (dSP_295_d[7:0] ), //i
    .b   (dSP_295_b[7:0] ), //i
    .p   (dSP_295_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_296 (
    .a   (dSP_296_a[7:0] ), //i
    .d   (dSP_296_d[7:0] ), //i
    .b   (dSP_296_b[7:0] ), //i
    .p   (dSP_296_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_297 (
    .a   (dSP_297_a[7:0] ), //i
    .d   (dSP_297_d[7:0] ), //i
    .b   (dSP_297_b[7:0] ), //i
    .p   (dSP_297_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_298 (
    .a   (dSP_298_a[7:0] ), //i
    .d   (dSP_298_d[7:0] ), //i
    .b   (dSP_298_b[7:0] ), //i
    .p   (dSP_298_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_299 (
    .a   (dSP_299_a[7:0] ), //i
    .d   (dSP_299_d[7:0] ), //i
    .b   (dSP_299_b[7:0] ), //i
    .p   (dSP_299_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_300 (
    .a   (dSP_300_a[7:0] ), //i
    .d   (dSP_300_d[7:0] ), //i
    .b   (dSP_300_b[7:0] ), //i
    .p   (dSP_300_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_301 (
    .a   (dSP_301_a[7:0] ), //i
    .d   (dSP_301_d[7:0] ), //i
    .b   (dSP_301_b[7:0] ), //i
    .p   (dSP_301_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_302 (
    .a   (dSP_302_a[7:0] ), //i
    .d   (dSP_302_d[7:0] ), //i
    .b   (dSP_302_b[7:0] ), //i
    .p   (dSP_302_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_303 (
    .a   (dSP_303_a[7:0] ), //i
    .d   (dSP_303_d[7:0] ), //i
    .b   (dSP_303_b[7:0] ), //i
    .p   (dSP_303_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_304 (
    .a   (dSP_304_a[7:0] ), //i
    .d   (dSP_304_d[7:0] ), //i
    .b   (dSP_304_b[7:0] ), //i
    .p   (dSP_304_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_305 (
    .a   (dSP_305_a[7:0] ), //i
    .d   (dSP_305_d[7:0] ), //i
    .b   (dSP_305_b[7:0] ), //i
    .p   (dSP_305_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_306 (
    .a   (dSP_306_a[7:0] ), //i
    .d   (dSP_306_d[7:0] ), //i
    .b   (dSP_306_b[7:0] ), //i
    .p   (dSP_306_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_307 (
    .a   (dSP_307_a[7:0] ), //i
    .d   (dSP_307_d[7:0] ), //i
    .b   (dSP_307_b[7:0] ), //i
    .p   (dSP_307_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_308 (
    .a   (dSP_308_a[7:0] ), //i
    .d   (dSP_308_d[7:0] ), //i
    .b   (dSP_308_b[7:0] ), //i
    .p   (dSP_308_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_309 (
    .a   (dSP_309_a[7:0] ), //i
    .d   (dSP_309_d[7:0] ), //i
    .b   (dSP_309_b[7:0] ), //i
    .p   (dSP_309_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_310 (
    .a   (dSP_310_a[7:0] ), //i
    .d   (dSP_310_d[7:0] ), //i
    .b   (dSP_310_b[7:0] ), //i
    .p   (dSP_310_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_311 (
    .a   (dSP_311_a[7:0] ), //i
    .d   (dSP_311_d[7:0] ), //i
    .b   (dSP_311_b[7:0] ), //i
    .p   (dSP_311_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_312 (
    .a   (dSP_312_a[7:0] ), //i
    .d   (dSP_312_d[7:0] ), //i
    .b   (dSP_312_b[7:0] ), //i
    .p   (dSP_312_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_313 (
    .a   (dSP_313_a[7:0] ), //i
    .d   (dSP_313_d[7:0] ), //i
    .b   (dSP_313_b[7:0] ), //i
    .p   (dSP_313_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_314 (
    .a   (dSP_314_a[7:0] ), //i
    .d   (dSP_314_d[7:0] ), //i
    .b   (dSP_314_b[7:0] ), //i
    .p   (dSP_314_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_315 (
    .a   (dSP_315_a[7:0] ), //i
    .d   (dSP_315_d[7:0] ), //i
    .b   (dSP_315_b[7:0] ), //i
    .p   (dSP_315_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_316 (
    .a   (dSP_316_a[7:0] ), //i
    .d   (dSP_316_d[7:0] ), //i
    .b   (dSP_316_b[7:0] ), //i
    .p   (dSP_316_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_317 (
    .a   (dSP_317_a[7:0] ), //i
    .d   (dSP_317_d[7:0] ), //i
    .b   (dSP_317_b[7:0] ), //i
    .p   (dSP_317_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_318 (
    .a   (dSP_318_a[7:0] ), //i
    .d   (dSP_318_d[7:0] ), //i
    .b   (dSP_318_b[7:0] ), //i
    .p   (dSP_318_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_319 (
    .a   (dSP_319_a[7:0] ), //i
    .d   (dSP_319_d[7:0] ), //i
    .b   (dSP_319_b[7:0] ), //i
    .p   (dSP_319_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_320 (
    .a   (dSP_320_a[7:0] ), //i
    .d   (dSP_320_d[7:0] ), //i
    .b   (dSP_320_b[7:0] ), //i
    .p   (dSP_320_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_321 (
    .a   (dSP_321_a[7:0] ), //i
    .d   (dSP_321_d[7:0] ), //i
    .b   (dSP_321_b[7:0] ), //i
    .p   (dSP_321_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_322 (
    .a   (dSP_322_a[7:0] ), //i
    .d   (dSP_322_d[7:0] ), //i
    .b   (dSP_322_b[7:0] ), //i
    .p   (dSP_322_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_323 (
    .a   (dSP_323_a[7:0] ), //i
    .d   (dSP_323_d[7:0] ), //i
    .b   (dSP_323_b[7:0] ), //i
    .p   (dSP_323_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_324 (
    .a   (dSP_324_a[7:0] ), //i
    .d   (dSP_324_d[7:0] ), //i
    .b   (dSP_324_b[7:0] ), //i
    .p   (dSP_324_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_325 (
    .a   (dSP_325_a[7:0] ), //i
    .d   (dSP_325_d[7:0] ), //i
    .b   (dSP_325_b[7:0] ), //i
    .p   (dSP_325_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_326 (
    .a   (dSP_326_a[7:0] ), //i
    .d   (dSP_326_d[7:0] ), //i
    .b   (dSP_326_b[7:0] ), //i
    .p   (dSP_326_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_327 (
    .a   (dSP_327_a[7:0] ), //i
    .d   (dSP_327_d[7:0] ), //i
    .b   (dSP_327_b[7:0] ), //i
    .p   (dSP_327_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_328 (
    .a   (dSP_328_a[7:0] ), //i
    .d   (dSP_328_d[7:0] ), //i
    .b   (dSP_328_b[7:0] ), //i
    .p   (dSP_328_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_329 (
    .a   (dSP_329_a[7:0] ), //i
    .d   (dSP_329_d[7:0] ), //i
    .b   (dSP_329_b[7:0] ), //i
    .p   (dSP_329_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_330 (
    .a   (dSP_330_a[7:0] ), //i
    .d   (dSP_330_d[7:0] ), //i
    .b   (dSP_330_b[7:0] ), //i
    .p   (dSP_330_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_331 (
    .a   (dSP_331_a[7:0] ), //i
    .d   (dSP_331_d[7:0] ), //i
    .b   (dSP_331_b[7:0] ), //i
    .p   (dSP_331_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_332 (
    .a   (dSP_332_a[7:0] ), //i
    .d   (dSP_332_d[7:0] ), //i
    .b   (dSP_332_b[7:0] ), //i
    .p   (dSP_332_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_333 (
    .a   (dSP_333_a[7:0] ), //i
    .d   (dSP_333_d[7:0] ), //i
    .b   (dSP_333_b[7:0] ), //i
    .p   (dSP_333_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_334 (
    .a   (dSP_334_a[7:0] ), //i
    .d   (dSP_334_d[7:0] ), //i
    .b   (dSP_334_b[7:0] ), //i
    .p   (dSP_334_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_335 (
    .a   (dSP_335_a[7:0] ), //i
    .d   (dSP_335_d[7:0] ), //i
    .b   (dSP_335_b[7:0] ), //i
    .p   (dSP_335_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_336 (
    .a   (dSP_336_a[7:0] ), //i
    .d   (dSP_336_d[7:0] ), //i
    .b   (dSP_336_b[7:0] ), //i
    .p   (dSP_336_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_337 (
    .a   (dSP_337_a[7:0] ), //i
    .d   (dSP_337_d[7:0] ), //i
    .b   (dSP_337_b[7:0] ), //i
    .p   (dSP_337_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_338 (
    .a   (dSP_338_a[7:0] ), //i
    .d   (dSP_338_d[7:0] ), //i
    .b   (dSP_338_b[7:0] ), //i
    .p   (dSP_338_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_339 (
    .a   (dSP_339_a[7:0] ), //i
    .d   (dSP_339_d[7:0] ), //i
    .b   (dSP_339_b[7:0] ), //i
    .p   (dSP_339_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_340 (
    .a   (dSP_340_a[7:0] ), //i
    .d   (dSP_340_d[7:0] ), //i
    .b   (dSP_340_b[7:0] ), //i
    .p   (dSP_340_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_341 (
    .a   (dSP_341_a[7:0] ), //i
    .d   (dSP_341_d[7:0] ), //i
    .b   (dSP_341_b[7:0] ), //i
    .p   (dSP_341_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_342 (
    .a   (dSP_342_a[7:0] ), //i
    .d   (dSP_342_d[7:0] ), //i
    .b   (dSP_342_b[7:0] ), //i
    .p   (dSP_342_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_343 (
    .a   (dSP_343_a[7:0] ), //i
    .d   (dSP_343_d[7:0] ), //i
    .b   (dSP_343_b[7:0] ), //i
    .p   (dSP_343_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_344 (
    .a   (dSP_344_a[7:0] ), //i
    .d   (dSP_344_d[7:0] ), //i
    .b   (dSP_344_b[7:0] ), //i
    .p   (dSP_344_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_345 (
    .a   (dSP_345_a[7:0] ), //i
    .d   (dSP_345_d[7:0] ), //i
    .b   (dSP_345_b[7:0] ), //i
    .p   (dSP_345_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_346 (
    .a   (dSP_346_a[7:0] ), //i
    .d   (dSP_346_d[7:0] ), //i
    .b   (dSP_346_b[7:0] ), //i
    .p   (dSP_346_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_347 (
    .a   (dSP_347_a[7:0] ), //i
    .d   (dSP_347_d[7:0] ), //i
    .b   (dSP_347_b[7:0] ), //i
    .p   (dSP_347_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_348 (
    .a   (dSP_348_a[7:0] ), //i
    .d   (dSP_348_d[7:0] ), //i
    .b   (dSP_348_b[7:0] ), //i
    .p   (dSP_348_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_349 (
    .a   (dSP_349_a[7:0] ), //i
    .d   (dSP_349_d[7:0] ), //i
    .b   (dSP_349_b[7:0] ), //i
    .p   (dSP_349_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_350 (
    .a   (dSP_350_a[7:0] ), //i
    .d   (dSP_350_d[7:0] ), //i
    .b   (dSP_350_b[7:0] ), //i
    .p   (dSP_350_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_351 (
    .a   (dSP_351_a[7:0] ), //i
    .d   (dSP_351_d[7:0] ), //i
    .b   (dSP_351_b[7:0] ), //i
    .p   (dSP_351_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_352 (
    .a   (dSP_352_a[7:0] ), //i
    .d   (dSP_352_d[7:0] ), //i
    .b   (dSP_352_b[7:0] ), //i
    .p   (dSP_352_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_353 (
    .a   (dSP_353_a[7:0] ), //i
    .d   (dSP_353_d[7:0] ), //i
    .b   (dSP_353_b[7:0] ), //i
    .p   (dSP_353_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_354 (
    .a   (dSP_354_a[7:0] ), //i
    .d   (dSP_354_d[7:0] ), //i
    .b   (dSP_354_b[7:0] ), //i
    .p   (dSP_354_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_355 (
    .a   (dSP_355_a[7:0] ), //i
    .d   (dSP_355_d[7:0] ), //i
    .b   (dSP_355_b[7:0] ), //i
    .p   (dSP_355_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_356 (
    .a   (dSP_356_a[7:0] ), //i
    .d   (dSP_356_d[7:0] ), //i
    .b   (dSP_356_b[7:0] ), //i
    .p   (dSP_356_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_357 (
    .a   (dSP_357_a[7:0] ), //i
    .d   (dSP_357_d[7:0] ), //i
    .b   (dSP_357_b[7:0] ), //i
    .p   (dSP_357_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_358 (
    .a   (dSP_358_a[7:0] ), //i
    .d   (dSP_358_d[7:0] ), //i
    .b   (dSP_358_b[7:0] ), //i
    .p   (dSP_358_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_359 (
    .a   (dSP_359_a[7:0] ), //i
    .d   (dSP_359_d[7:0] ), //i
    .b   (dSP_359_b[7:0] ), //i
    .p   (dSP_359_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_360 (
    .a   (dSP_360_a[7:0] ), //i
    .d   (dSP_360_d[7:0] ), //i
    .b   (dSP_360_b[7:0] ), //i
    .p   (dSP_360_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_361 (
    .a   (dSP_361_a[7:0] ), //i
    .d   (dSP_361_d[7:0] ), //i
    .b   (dSP_361_b[7:0] ), //i
    .p   (dSP_361_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_362 (
    .a   (dSP_362_a[7:0] ), //i
    .d   (dSP_362_d[7:0] ), //i
    .b   (dSP_362_b[7:0] ), //i
    .p   (dSP_362_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_363 (
    .a   (dSP_363_a[7:0] ), //i
    .d   (dSP_363_d[7:0] ), //i
    .b   (dSP_363_b[7:0] ), //i
    .p   (dSP_363_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_364 (
    .a   (dSP_364_a[7:0] ), //i
    .d   (dSP_364_d[7:0] ), //i
    .b   (dSP_364_b[7:0] ), //i
    .p   (dSP_364_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_365 (
    .a   (dSP_365_a[7:0] ), //i
    .d   (dSP_365_d[7:0] ), //i
    .b   (dSP_365_b[7:0] ), //i
    .p   (dSP_365_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_366 (
    .a   (dSP_366_a[7:0] ), //i
    .d   (dSP_366_d[7:0] ), //i
    .b   (dSP_366_b[7:0] ), //i
    .p   (dSP_366_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_367 (
    .a   (dSP_367_a[7:0] ), //i
    .d   (dSP_367_d[7:0] ), //i
    .b   (dSP_367_b[7:0] ), //i
    .p   (dSP_367_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_368 (
    .a   (dSP_368_a[7:0] ), //i
    .d   (dSP_368_d[7:0] ), //i
    .b   (dSP_368_b[7:0] ), //i
    .p   (dSP_368_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_369 (
    .a   (dSP_369_a[7:0] ), //i
    .d   (dSP_369_d[7:0] ), //i
    .b   (dSP_369_b[7:0] ), //i
    .p   (dSP_369_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_370 (
    .a   (dSP_370_a[7:0] ), //i
    .d   (dSP_370_d[7:0] ), //i
    .b   (dSP_370_b[7:0] ), //i
    .p   (dSP_370_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_371 (
    .a   (dSP_371_a[7:0] ), //i
    .d   (dSP_371_d[7:0] ), //i
    .b   (dSP_371_b[7:0] ), //i
    .p   (dSP_371_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_372 (
    .a   (dSP_372_a[7:0] ), //i
    .d   (dSP_372_d[7:0] ), //i
    .b   (dSP_372_b[7:0] ), //i
    .p   (dSP_372_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_373 (
    .a   (dSP_373_a[7:0] ), //i
    .d   (dSP_373_d[7:0] ), //i
    .b   (dSP_373_b[7:0] ), //i
    .p   (dSP_373_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_374 (
    .a   (dSP_374_a[7:0] ), //i
    .d   (dSP_374_d[7:0] ), //i
    .b   (dSP_374_b[7:0] ), //i
    .p   (dSP_374_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_375 (
    .a   (dSP_375_a[7:0] ), //i
    .d   (dSP_375_d[7:0] ), //i
    .b   (dSP_375_b[7:0] ), //i
    .p   (dSP_375_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_376 (
    .a   (dSP_376_a[7:0] ), //i
    .d   (dSP_376_d[7:0] ), //i
    .b   (dSP_376_b[7:0] ), //i
    .p   (dSP_376_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_377 (
    .a   (dSP_377_a[7:0] ), //i
    .d   (dSP_377_d[7:0] ), //i
    .b   (dSP_377_b[7:0] ), //i
    .p   (dSP_377_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_378 (
    .a   (dSP_378_a[7:0] ), //i
    .d   (dSP_378_d[7:0] ), //i
    .b   (dSP_378_b[7:0] ), //i
    .p   (dSP_378_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_379 (
    .a   (dSP_379_a[7:0] ), //i
    .d   (dSP_379_d[7:0] ), //i
    .b   (dSP_379_b[7:0] ), //i
    .p   (dSP_379_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_380 (
    .a   (dSP_380_a[7:0] ), //i
    .d   (dSP_380_d[7:0] ), //i
    .b   (dSP_380_b[7:0] ), //i
    .p   (dSP_380_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_381 (
    .a   (dSP_381_a[7:0] ), //i
    .d   (dSP_381_d[7:0] ), //i
    .b   (dSP_381_b[7:0] ), //i
    .p   (dSP_381_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_382 (
    .a   (dSP_382_a[7:0] ), //i
    .d   (dSP_382_d[7:0] ), //i
    .b   (dSP_382_b[7:0] ), //i
    .p   (dSP_382_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_383 (
    .a   (dSP_383_a[7:0] ), //i
    .d   (dSP_383_d[7:0] ), //i
    .b   (dSP_383_b[7:0] ), //i
    .p   (dSP_383_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_384 (
    .a   (dSP_384_a[7:0] ), //i
    .d   (dSP_384_d[7:0] ), //i
    .b   (dSP_384_b[7:0] ), //i
    .p   (dSP_384_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_385 (
    .a   (dSP_385_a[7:0] ), //i
    .d   (dSP_385_d[7:0] ), //i
    .b   (dSP_385_b[7:0] ), //i
    .p   (dSP_385_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_386 (
    .a   (dSP_386_a[7:0] ), //i
    .d   (dSP_386_d[7:0] ), //i
    .b   (dSP_386_b[7:0] ), //i
    .p   (dSP_386_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_387 (
    .a   (dSP_387_a[7:0] ), //i
    .d   (dSP_387_d[7:0] ), //i
    .b   (dSP_387_b[7:0] ), //i
    .p   (dSP_387_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_388 (
    .a   (dSP_388_a[7:0] ), //i
    .d   (dSP_388_d[7:0] ), //i
    .b   (dSP_388_b[7:0] ), //i
    .p   (dSP_388_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_389 (
    .a   (dSP_389_a[7:0] ), //i
    .d   (dSP_389_d[7:0] ), //i
    .b   (dSP_389_b[7:0] ), //i
    .p   (dSP_389_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_390 (
    .a   (dSP_390_a[7:0] ), //i
    .d   (dSP_390_d[7:0] ), //i
    .b   (dSP_390_b[7:0] ), //i
    .p   (dSP_390_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_391 (
    .a   (dSP_391_a[7:0] ), //i
    .d   (dSP_391_d[7:0] ), //i
    .b   (dSP_391_b[7:0] ), //i
    .p   (dSP_391_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_392 (
    .a   (dSP_392_a[7:0] ), //i
    .d   (dSP_392_d[7:0] ), //i
    .b   (dSP_392_b[7:0] ), //i
    .p   (dSP_392_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_393 (
    .a   (dSP_393_a[7:0] ), //i
    .d   (dSP_393_d[7:0] ), //i
    .b   (dSP_393_b[7:0] ), //i
    .p   (dSP_393_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_394 (
    .a   (dSP_394_a[7:0] ), //i
    .d   (dSP_394_d[7:0] ), //i
    .b   (dSP_394_b[7:0] ), //i
    .p   (dSP_394_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_395 (
    .a   (dSP_395_a[7:0] ), //i
    .d   (dSP_395_d[7:0] ), //i
    .b   (dSP_395_b[7:0] ), //i
    .p   (dSP_395_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_396 (
    .a   (dSP_396_a[7:0] ), //i
    .d   (dSP_396_d[7:0] ), //i
    .b   (dSP_396_b[7:0] ), //i
    .p   (dSP_396_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_397 (
    .a   (dSP_397_a[7:0] ), //i
    .d   (dSP_397_d[7:0] ), //i
    .b   (dSP_397_b[7:0] ), //i
    .p   (dSP_397_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_398 (
    .a   (dSP_398_a[7:0] ), //i
    .d   (dSP_398_d[7:0] ), //i
    .b   (dSP_398_b[7:0] ), //i
    .p   (dSP_398_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_399 (
    .a   (dSP_399_a[7:0] ), //i
    .d   (dSP_399_d[7:0] ), //i
    .b   (dSP_399_b[7:0] ), //i
    .p   (dSP_399_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_400 (
    .a   (dSP_400_a[7:0] ), //i
    .d   (dSP_400_d[7:0] ), //i
    .b   (dSP_400_b[7:0] ), //i
    .p   (dSP_400_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_401 (
    .a   (dSP_401_a[7:0] ), //i
    .d   (dSP_401_d[7:0] ), //i
    .b   (dSP_401_b[7:0] ), //i
    .p   (dSP_401_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_402 (
    .a   (dSP_402_a[7:0] ), //i
    .d   (dSP_402_d[7:0] ), //i
    .b   (dSP_402_b[7:0] ), //i
    .p   (dSP_402_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_403 (
    .a   (dSP_403_a[7:0] ), //i
    .d   (dSP_403_d[7:0] ), //i
    .b   (dSP_403_b[7:0] ), //i
    .p   (dSP_403_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_404 (
    .a   (dSP_404_a[7:0] ), //i
    .d   (dSP_404_d[7:0] ), //i
    .b   (dSP_404_b[7:0] ), //i
    .p   (dSP_404_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_405 (
    .a   (dSP_405_a[7:0] ), //i
    .d   (dSP_405_d[7:0] ), //i
    .b   (dSP_405_b[7:0] ), //i
    .p   (dSP_405_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_406 (
    .a   (dSP_406_a[7:0] ), //i
    .d   (dSP_406_d[7:0] ), //i
    .b   (dSP_406_b[7:0] ), //i
    .p   (dSP_406_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_407 (
    .a   (dSP_407_a[7:0] ), //i
    .d   (dSP_407_d[7:0] ), //i
    .b   (dSP_407_b[7:0] ), //i
    .p   (dSP_407_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_408 (
    .a   (dSP_408_a[7:0] ), //i
    .d   (dSP_408_d[7:0] ), //i
    .b   (dSP_408_b[7:0] ), //i
    .p   (dSP_408_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_409 (
    .a   (dSP_409_a[7:0] ), //i
    .d   (dSP_409_d[7:0] ), //i
    .b   (dSP_409_b[7:0] ), //i
    .p   (dSP_409_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_410 (
    .a   (dSP_410_a[7:0] ), //i
    .d   (dSP_410_d[7:0] ), //i
    .b   (dSP_410_b[7:0] ), //i
    .p   (dSP_410_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_411 (
    .a   (dSP_411_a[7:0] ), //i
    .d   (dSP_411_d[7:0] ), //i
    .b   (dSP_411_b[7:0] ), //i
    .p   (dSP_411_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_412 (
    .a   (dSP_412_a[7:0] ), //i
    .d   (dSP_412_d[7:0] ), //i
    .b   (dSP_412_b[7:0] ), //i
    .p   (dSP_412_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_413 (
    .a   (dSP_413_a[7:0] ), //i
    .d   (dSP_413_d[7:0] ), //i
    .b   (dSP_413_b[7:0] ), //i
    .p   (dSP_413_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_414 (
    .a   (dSP_414_a[7:0] ), //i
    .d   (dSP_414_d[7:0] ), //i
    .b   (dSP_414_b[7:0] ), //i
    .p   (dSP_414_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_415 (
    .a   (dSP_415_a[7:0] ), //i
    .d   (dSP_415_d[7:0] ), //i
    .b   (dSP_415_b[7:0] ), //i
    .p   (dSP_415_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_416 (
    .a   (dSP_416_a[7:0] ), //i
    .d   (dSP_416_d[7:0] ), //i
    .b   (dSP_416_b[7:0] ), //i
    .p   (dSP_416_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_417 (
    .a   (dSP_417_a[7:0] ), //i
    .d   (dSP_417_d[7:0] ), //i
    .b   (dSP_417_b[7:0] ), //i
    .p   (dSP_417_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_418 (
    .a   (dSP_418_a[7:0] ), //i
    .d   (dSP_418_d[7:0] ), //i
    .b   (dSP_418_b[7:0] ), //i
    .p   (dSP_418_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_419 (
    .a   (dSP_419_a[7:0] ), //i
    .d   (dSP_419_d[7:0] ), //i
    .b   (dSP_419_b[7:0] ), //i
    .p   (dSP_419_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_420 (
    .a   (dSP_420_a[7:0] ), //i
    .d   (dSP_420_d[7:0] ), //i
    .b   (dSP_420_b[7:0] ), //i
    .p   (dSP_420_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_421 (
    .a   (dSP_421_a[7:0] ), //i
    .d   (dSP_421_d[7:0] ), //i
    .b   (dSP_421_b[7:0] ), //i
    .p   (dSP_421_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_422 (
    .a   (dSP_422_a[7:0] ), //i
    .d   (dSP_422_d[7:0] ), //i
    .b   (dSP_422_b[7:0] ), //i
    .p   (dSP_422_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_423 (
    .a   (dSP_423_a[7:0] ), //i
    .d   (dSP_423_d[7:0] ), //i
    .b   (dSP_423_b[7:0] ), //i
    .p   (dSP_423_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_424 (
    .a   (dSP_424_a[7:0] ), //i
    .d   (dSP_424_d[7:0] ), //i
    .b   (dSP_424_b[7:0] ), //i
    .p   (dSP_424_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_425 (
    .a   (dSP_425_a[7:0] ), //i
    .d   (dSP_425_d[7:0] ), //i
    .b   (dSP_425_b[7:0] ), //i
    .p   (dSP_425_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_426 (
    .a   (dSP_426_a[7:0] ), //i
    .d   (dSP_426_d[7:0] ), //i
    .b   (dSP_426_b[7:0] ), //i
    .p   (dSP_426_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_427 (
    .a   (dSP_427_a[7:0] ), //i
    .d   (dSP_427_d[7:0] ), //i
    .b   (dSP_427_b[7:0] ), //i
    .p   (dSP_427_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_428 (
    .a   (dSP_428_a[7:0] ), //i
    .d   (dSP_428_d[7:0] ), //i
    .b   (dSP_428_b[7:0] ), //i
    .p   (dSP_428_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_429 (
    .a   (dSP_429_a[7:0] ), //i
    .d   (dSP_429_d[7:0] ), //i
    .b   (dSP_429_b[7:0] ), //i
    .p   (dSP_429_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_430 (
    .a   (dSP_430_a[7:0] ), //i
    .d   (dSP_430_d[7:0] ), //i
    .b   (dSP_430_b[7:0] ), //i
    .p   (dSP_430_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_431 (
    .a   (dSP_431_a[7:0] ), //i
    .d   (dSP_431_d[7:0] ), //i
    .b   (dSP_431_b[7:0] ), //i
    .p   (dSP_431_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_432 (
    .a   (dSP_432_a[7:0] ), //i
    .d   (dSP_432_d[7:0] ), //i
    .b   (dSP_432_b[7:0] ), //i
    .p   (dSP_432_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_433 (
    .a   (dSP_433_a[7:0] ), //i
    .d   (dSP_433_d[7:0] ), //i
    .b   (dSP_433_b[7:0] ), //i
    .p   (dSP_433_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_434 (
    .a   (dSP_434_a[7:0] ), //i
    .d   (dSP_434_d[7:0] ), //i
    .b   (dSP_434_b[7:0] ), //i
    .p   (dSP_434_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_435 (
    .a   (dSP_435_a[7:0] ), //i
    .d   (dSP_435_d[7:0] ), //i
    .b   (dSP_435_b[7:0] ), //i
    .p   (dSP_435_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_436 (
    .a   (dSP_436_a[7:0] ), //i
    .d   (dSP_436_d[7:0] ), //i
    .b   (dSP_436_b[7:0] ), //i
    .p   (dSP_436_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_437 (
    .a   (dSP_437_a[7:0] ), //i
    .d   (dSP_437_d[7:0] ), //i
    .b   (dSP_437_b[7:0] ), //i
    .p   (dSP_437_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_438 (
    .a   (dSP_438_a[7:0] ), //i
    .d   (dSP_438_d[7:0] ), //i
    .b   (dSP_438_b[7:0] ), //i
    .p   (dSP_438_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_439 (
    .a   (dSP_439_a[7:0] ), //i
    .d   (dSP_439_d[7:0] ), //i
    .b   (dSP_439_b[7:0] ), //i
    .p   (dSP_439_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_440 (
    .a   (dSP_440_a[7:0] ), //i
    .d   (dSP_440_d[7:0] ), //i
    .b   (dSP_440_b[7:0] ), //i
    .p   (dSP_440_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_441 (
    .a   (dSP_441_a[7:0] ), //i
    .d   (dSP_441_d[7:0] ), //i
    .b   (dSP_441_b[7:0] ), //i
    .p   (dSP_441_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_442 (
    .a   (dSP_442_a[7:0] ), //i
    .d   (dSP_442_d[7:0] ), //i
    .b   (dSP_442_b[7:0] ), //i
    .p   (dSP_442_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_443 (
    .a   (dSP_443_a[7:0] ), //i
    .d   (dSP_443_d[7:0] ), //i
    .b   (dSP_443_b[7:0] ), //i
    .p   (dSP_443_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_444 (
    .a   (dSP_444_a[7:0] ), //i
    .d   (dSP_444_d[7:0] ), //i
    .b   (dSP_444_b[7:0] ), //i
    .p   (dSP_444_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_445 (
    .a   (dSP_445_a[7:0] ), //i
    .d   (dSP_445_d[7:0] ), //i
    .b   (dSP_445_b[7:0] ), //i
    .p   (dSP_445_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_446 (
    .a   (dSP_446_a[7:0] ), //i
    .d   (dSP_446_d[7:0] ), //i
    .b   (dSP_446_b[7:0] ), //i
    .p   (dSP_446_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_447 (
    .a   (dSP_447_a[7:0] ), //i
    .d   (dSP_447_d[7:0] ), //i
    .b   (dSP_447_b[7:0] ), //i
    .p   (dSP_447_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_448 (
    .a   (dSP_448_a[7:0] ), //i
    .d   (dSP_448_d[7:0] ), //i
    .b   (dSP_448_b[7:0] ), //i
    .p   (dSP_448_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_449 (
    .a   (dSP_449_a[7:0] ), //i
    .d   (dSP_449_d[7:0] ), //i
    .b   (dSP_449_b[7:0] ), //i
    .p   (dSP_449_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_450 (
    .a   (dSP_450_a[7:0] ), //i
    .d   (dSP_450_d[7:0] ), //i
    .b   (dSP_450_b[7:0] ), //i
    .p   (dSP_450_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_451 (
    .a   (dSP_451_a[7:0] ), //i
    .d   (dSP_451_d[7:0] ), //i
    .b   (dSP_451_b[7:0] ), //i
    .p   (dSP_451_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_452 (
    .a   (dSP_452_a[7:0] ), //i
    .d   (dSP_452_d[7:0] ), //i
    .b   (dSP_452_b[7:0] ), //i
    .p   (dSP_452_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_453 (
    .a   (dSP_453_a[7:0] ), //i
    .d   (dSP_453_d[7:0] ), //i
    .b   (dSP_453_b[7:0] ), //i
    .p   (dSP_453_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_454 (
    .a   (dSP_454_a[7:0] ), //i
    .d   (dSP_454_d[7:0] ), //i
    .b   (dSP_454_b[7:0] ), //i
    .p   (dSP_454_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_455 (
    .a   (dSP_455_a[7:0] ), //i
    .d   (dSP_455_d[7:0] ), //i
    .b   (dSP_455_b[7:0] ), //i
    .p   (dSP_455_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_456 (
    .a   (dSP_456_a[7:0] ), //i
    .d   (dSP_456_d[7:0] ), //i
    .b   (dSP_456_b[7:0] ), //i
    .p   (dSP_456_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_457 (
    .a   (dSP_457_a[7:0] ), //i
    .d   (dSP_457_d[7:0] ), //i
    .b   (dSP_457_b[7:0] ), //i
    .p   (dSP_457_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_458 (
    .a   (dSP_458_a[7:0] ), //i
    .d   (dSP_458_d[7:0] ), //i
    .b   (dSP_458_b[7:0] ), //i
    .p   (dSP_458_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_459 (
    .a   (dSP_459_a[7:0] ), //i
    .d   (dSP_459_d[7:0] ), //i
    .b   (dSP_459_b[7:0] ), //i
    .p   (dSP_459_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_460 (
    .a   (dSP_460_a[7:0] ), //i
    .d   (dSP_460_d[7:0] ), //i
    .b   (dSP_460_b[7:0] ), //i
    .p   (dSP_460_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_461 (
    .a   (dSP_461_a[7:0] ), //i
    .d   (dSP_461_d[7:0] ), //i
    .b   (dSP_461_b[7:0] ), //i
    .p   (dSP_461_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_462 (
    .a   (dSP_462_a[7:0] ), //i
    .d   (dSP_462_d[7:0] ), //i
    .b   (dSP_462_b[7:0] ), //i
    .p   (dSP_462_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_463 (
    .a   (dSP_463_a[7:0] ), //i
    .d   (dSP_463_d[7:0] ), //i
    .b   (dSP_463_b[7:0] ), //i
    .p   (dSP_463_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_464 (
    .a   (dSP_464_a[7:0] ), //i
    .d   (dSP_464_d[7:0] ), //i
    .b   (dSP_464_b[7:0] ), //i
    .p   (dSP_464_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_465 (
    .a   (dSP_465_a[7:0] ), //i
    .d   (dSP_465_d[7:0] ), //i
    .b   (dSP_465_b[7:0] ), //i
    .p   (dSP_465_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_466 (
    .a   (dSP_466_a[7:0] ), //i
    .d   (dSP_466_d[7:0] ), //i
    .b   (dSP_466_b[7:0] ), //i
    .p   (dSP_466_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_467 (
    .a   (dSP_467_a[7:0] ), //i
    .d   (dSP_467_d[7:0] ), //i
    .b   (dSP_467_b[7:0] ), //i
    .p   (dSP_467_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_468 (
    .a   (dSP_468_a[7:0] ), //i
    .d   (dSP_468_d[7:0] ), //i
    .b   (dSP_468_b[7:0] ), //i
    .p   (dSP_468_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_469 (
    .a   (dSP_469_a[7:0] ), //i
    .d   (dSP_469_d[7:0] ), //i
    .b   (dSP_469_b[7:0] ), //i
    .p   (dSP_469_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_470 (
    .a   (dSP_470_a[7:0] ), //i
    .d   (dSP_470_d[7:0] ), //i
    .b   (dSP_470_b[7:0] ), //i
    .p   (dSP_470_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_471 (
    .a   (dSP_471_a[7:0] ), //i
    .d   (dSP_471_d[7:0] ), //i
    .b   (dSP_471_b[7:0] ), //i
    .p   (dSP_471_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_472 (
    .a   (dSP_472_a[7:0] ), //i
    .d   (dSP_472_d[7:0] ), //i
    .b   (dSP_472_b[7:0] ), //i
    .p   (dSP_472_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_473 (
    .a   (dSP_473_a[7:0] ), //i
    .d   (dSP_473_d[7:0] ), //i
    .b   (dSP_473_b[7:0] ), //i
    .p   (dSP_473_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_474 (
    .a   (dSP_474_a[7:0] ), //i
    .d   (dSP_474_d[7:0] ), //i
    .b   (dSP_474_b[7:0] ), //i
    .p   (dSP_474_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_475 (
    .a   (dSP_475_a[7:0] ), //i
    .d   (dSP_475_d[7:0] ), //i
    .b   (dSP_475_b[7:0] ), //i
    .p   (dSP_475_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_476 (
    .a   (dSP_476_a[7:0] ), //i
    .d   (dSP_476_d[7:0] ), //i
    .b   (dSP_476_b[7:0] ), //i
    .p   (dSP_476_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_477 (
    .a   (dSP_477_a[7:0] ), //i
    .d   (dSP_477_d[7:0] ), //i
    .b   (dSP_477_b[7:0] ), //i
    .p   (dSP_477_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_478 (
    .a   (dSP_478_a[7:0] ), //i
    .d   (dSP_478_d[7:0] ), //i
    .b   (dSP_478_b[7:0] ), //i
    .p   (dSP_478_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_479 (
    .a   (dSP_479_a[7:0] ), //i
    .d   (dSP_479_d[7:0] ), //i
    .b   (dSP_479_b[7:0] ), //i
    .p   (dSP_479_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_480 (
    .a   (dSP_480_a[7:0] ), //i
    .d   (dSP_480_d[7:0] ), //i
    .b   (dSP_480_b[7:0] ), //i
    .p   (dSP_480_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_481 (
    .a   (dSP_481_a[7:0] ), //i
    .d   (dSP_481_d[7:0] ), //i
    .b   (dSP_481_b[7:0] ), //i
    .p   (dSP_481_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_482 (
    .a   (dSP_482_a[7:0] ), //i
    .d   (dSP_482_d[7:0] ), //i
    .b   (dSP_482_b[7:0] ), //i
    .p   (dSP_482_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_483 (
    .a   (dSP_483_a[7:0] ), //i
    .d   (dSP_483_d[7:0] ), //i
    .b   (dSP_483_b[7:0] ), //i
    .p   (dSP_483_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_484 (
    .a   (dSP_484_a[7:0] ), //i
    .d   (dSP_484_d[7:0] ), //i
    .b   (dSP_484_b[7:0] ), //i
    .p   (dSP_484_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_485 (
    .a   (dSP_485_a[7:0] ), //i
    .d   (dSP_485_d[7:0] ), //i
    .b   (dSP_485_b[7:0] ), //i
    .p   (dSP_485_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_486 (
    .a   (dSP_486_a[7:0] ), //i
    .d   (dSP_486_d[7:0] ), //i
    .b   (dSP_486_b[7:0] ), //i
    .p   (dSP_486_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_487 (
    .a   (dSP_487_a[7:0] ), //i
    .d   (dSP_487_d[7:0] ), //i
    .b   (dSP_487_b[7:0] ), //i
    .p   (dSP_487_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_488 (
    .a   (dSP_488_a[7:0] ), //i
    .d   (dSP_488_d[7:0] ), //i
    .b   (dSP_488_b[7:0] ), //i
    .p   (dSP_488_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_489 (
    .a   (dSP_489_a[7:0] ), //i
    .d   (dSP_489_d[7:0] ), //i
    .b   (dSP_489_b[7:0] ), //i
    .p   (dSP_489_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_490 (
    .a   (dSP_490_a[7:0] ), //i
    .d   (dSP_490_d[7:0] ), //i
    .b   (dSP_490_b[7:0] ), //i
    .p   (dSP_490_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_491 (
    .a   (dSP_491_a[7:0] ), //i
    .d   (dSP_491_d[7:0] ), //i
    .b   (dSP_491_b[7:0] ), //i
    .p   (dSP_491_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_492 (
    .a   (dSP_492_a[7:0] ), //i
    .d   (dSP_492_d[7:0] ), //i
    .b   (dSP_492_b[7:0] ), //i
    .p   (dSP_492_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_493 (
    .a   (dSP_493_a[7:0] ), //i
    .d   (dSP_493_d[7:0] ), //i
    .b   (dSP_493_b[7:0] ), //i
    .p   (dSP_493_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_494 (
    .a   (dSP_494_a[7:0] ), //i
    .d   (dSP_494_d[7:0] ), //i
    .b   (dSP_494_b[7:0] ), //i
    .p   (dSP_494_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_495 (
    .a   (dSP_495_a[7:0] ), //i
    .d   (dSP_495_d[7:0] ), //i
    .b   (dSP_495_b[7:0] ), //i
    .p   (dSP_495_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_496 (
    .a   (dSP_496_a[7:0] ), //i
    .d   (dSP_496_d[7:0] ), //i
    .b   (dSP_496_b[7:0] ), //i
    .p   (dSP_496_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_497 (
    .a   (dSP_497_a[7:0] ), //i
    .d   (dSP_497_d[7:0] ), //i
    .b   (dSP_497_b[7:0] ), //i
    .p   (dSP_497_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_498 (
    .a   (dSP_498_a[7:0] ), //i
    .d   (dSP_498_d[7:0] ), //i
    .b   (dSP_498_b[7:0] ), //i
    .p   (dSP_498_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_499 (
    .a   (dSP_499_a[7:0] ), //i
    .d   (dSP_499_d[7:0] ), //i
    .b   (dSP_499_b[7:0] ), //i
    .p   (dSP_499_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_500 (
    .a   (dSP_500_a[7:0] ), //i
    .d   (dSP_500_d[7:0] ), //i
    .b   (dSP_500_b[7:0] ), //i
    .p   (dSP_500_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_501 (
    .a   (dSP_501_a[7:0] ), //i
    .d   (dSP_501_d[7:0] ), //i
    .b   (dSP_501_b[7:0] ), //i
    .p   (dSP_501_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_502 (
    .a   (dSP_502_a[7:0] ), //i
    .d   (dSP_502_d[7:0] ), //i
    .b   (dSP_502_b[7:0] ), //i
    .p   (dSP_502_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_503 (
    .a   (dSP_503_a[7:0] ), //i
    .d   (dSP_503_d[7:0] ), //i
    .b   (dSP_503_b[7:0] ), //i
    .p   (dSP_503_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_504 (
    .a   (dSP_504_a[7:0] ), //i
    .d   (dSP_504_d[7:0] ), //i
    .b   (dSP_504_b[7:0] ), //i
    .p   (dSP_504_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_505 (
    .a   (dSP_505_a[7:0] ), //i
    .d   (dSP_505_d[7:0] ), //i
    .b   (dSP_505_b[7:0] ), //i
    .p   (dSP_505_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_506 (
    .a   (dSP_506_a[7:0] ), //i
    .d   (dSP_506_d[7:0] ), //i
    .b   (dSP_506_b[7:0] ), //i
    .p   (dSP_506_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_507 (
    .a   (dSP_507_a[7:0] ), //i
    .d   (dSP_507_d[7:0] ), //i
    .b   (dSP_507_b[7:0] ), //i
    .p   (dSP_507_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_508 (
    .a   (dSP_508_a[7:0] ), //i
    .d   (dSP_508_d[7:0] ), //i
    .b   (dSP_508_b[7:0] ), //i
    .p   (dSP_508_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_509 (
    .a   (dSP_509_a[7:0] ), //i
    .d   (dSP_509_d[7:0] ), //i
    .b   (dSP_509_b[7:0] ), //i
    .p   (dSP_509_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_510 (
    .a   (dSP_510_a[7:0] ), //i
    .d   (dSP_510_d[7:0] ), //i
    .b   (dSP_510_b[7:0] ), //i
    .p   (dSP_510_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_511 (
    .a   (dSP_511_a[7:0] ), //i
    .d   (dSP_511_d[7:0] ), //i
    .b   (dSP_511_b[7:0] ), //i
    .p   (dSP_511_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_512 (
    .a   (dSP_512_a[7:0] ), //i
    .d   (dSP_512_d[7:0] ), //i
    .b   (dSP_512_b[7:0] ), //i
    .p   (dSP_512_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_513 (
    .a   (dSP_513_a[7:0] ), //i
    .d   (dSP_513_d[7:0] ), //i
    .b   (dSP_513_b[7:0] ), //i
    .p   (dSP_513_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_514 (
    .a   (dSP_514_a[7:0] ), //i
    .d   (dSP_514_d[7:0] ), //i
    .b   (dSP_514_b[7:0] ), //i
    .p   (dSP_514_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_515 (
    .a   (dSP_515_a[7:0] ), //i
    .d   (dSP_515_d[7:0] ), //i
    .b   (dSP_515_b[7:0] ), //i
    .p   (dSP_515_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_516 (
    .a   (dSP_516_a[7:0] ), //i
    .d   (dSP_516_d[7:0] ), //i
    .b   (dSP_516_b[7:0] ), //i
    .p   (dSP_516_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_517 (
    .a   (dSP_517_a[7:0] ), //i
    .d   (dSP_517_d[7:0] ), //i
    .b   (dSP_517_b[7:0] ), //i
    .p   (dSP_517_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_518 (
    .a   (dSP_518_a[7:0] ), //i
    .d   (dSP_518_d[7:0] ), //i
    .b   (dSP_518_b[7:0] ), //i
    .p   (dSP_518_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_519 (
    .a   (dSP_519_a[7:0] ), //i
    .d   (dSP_519_d[7:0] ), //i
    .b   (dSP_519_b[7:0] ), //i
    .p   (dSP_519_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_520 (
    .a   (dSP_520_a[7:0] ), //i
    .d   (dSP_520_d[7:0] ), //i
    .b   (dSP_520_b[7:0] ), //i
    .p   (dSP_520_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_521 (
    .a   (dSP_521_a[7:0] ), //i
    .d   (dSP_521_d[7:0] ), //i
    .b   (dSP_521_b[7:0] ), //i
    .p   (dSP_521_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_522 (
    .a   (dSP_522_a[7:0] ), //i
    .d   (dSP_522_d[7:0] ), //i
    .b   (dSP_522_b[7:0] ), //i
    .p   (dSP_522_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_523 (
    .a   (dSP_523_a[7:0] ), //i
    .d   (dSP_523_d[7:0] ), //i
    .b   (dSP_523_b[7:0] ), //i
    .p   (dSP_523_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_524 (
    .a   (dSP_524_a[7:0] ), //i
    .d   (dSP_524_d[7:0] ), //i
    .b   (dSP_524_b[7:0] ), //i
    .p   (dSP_524_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_525 (
    .a   (dSP_525_a[7:0] ), //i
    .d   (dSP_525_d[7:0] ), //i
    .b   (dSP_525_b[7:0] ), //i
    .p   (dSP_525_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_526 (
    .a   (dSP_526_a[7:0] ), //i
    .d   (dSP_526_d[7:0] ), //i
    .b   (dSP_526_b[7:0] ), //i
    .p   (dSP_526_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_527 (
    .a   (dSP_527_a[7:0] ), //i
    .d   (dSP_527_d[7:0] ), //i
    .b   (dSP_527_b[7:0] ), //i
    .p   (dSP_527_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_528 (
    .a   (dSP_528_a[7:0] ), //i
    .d   (dSP_528_d[7:0] ), //i
    .b   (dSP_528_b[7:0] ), //i
    .p   (dSP_528_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_529 (
    .a   (dSP_529_a[7:0] ), //i
    .d   (dSP_529_d[7:0] ), //i
    .b   (dSP_529_b[7:0] ), //i
    .p   (dSP_529_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_530 (
    .a   (dSP_530_a[7:0] ), //i
    .d   (dSP_530_d[7:0] ), //i
    .b   (dSP_530_b[7:0] ), //i
    .p   (dSP_530_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_531 (
    .a   (dSP_531_a[7:0] ), //i
    .d   (dSP_531_d[7:0] ), //i
    .b   (dSP_531_b[7:0] ), //i
    .p   (dSP_531_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_532 (
    .a   (dSP_532_a[7:0] ), //i
    .d   (dSP_532_d[7:0] ), //i
    .b   (dSP_532_b[7:0] ), //i
    .p   (dSP_532_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_533 (
    .a   (dSP_533_a[7:0] ), //i
    .d   (dSP_533_d[7:0] ), //i
    .b   (dSP_533_b[7:0] ), //i
    .p   (dSP_533_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_534 (
    .a   (dSP_534_a[7:0] ), //i
    .d   (dSP_534_d[7:0] ), //i
    .b   (dSP_534_b[7:0] ), //i
    .p   (dSP_534_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_535 (
    .a   (dSP_535_a[7:0] ), //i
    .d   (dSP_535_d[7:0] ), //i
    .b   (dSP_535_b[7:0] ), //i
    .p   (dSP_535_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_536 (
    .a   (dSP_536_a[7:0] ), //i
    .d   (dSP_536_d[7:0] ), //i
    .b   (dSP_536_b[7:0] ), //i
    .p   (dSP_536_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_537 (
    .a   (dSP_537_a[7:0] ), //i
    .d   (dSP_537_d[7:0] ), //i
    .b   (dSP_537_b[7:0] ), //i
    .p   (dSP_537_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_538 (
    .a   (dSP_538_a[7:0] ), //i
    .d   (dSP_538_d[7:0] ), //i
    .b   (dSP_538_b[7:0] ), //i
    .p   (dSP_538_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_539 (
    .a   (dSP_539_a[7:0] ), //i
    .d   (dSP_539_d[7:0] ), //i
    .b   (dSP_539_b[7:0] ), //i
    .p   (dSP_539_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_540 (
    .a   (dSP_540_a[7:0] ), //i
    .d   (dSP_540_d[7:0] ), //i
    .b   (dSP_540_b[7:0] ), //i
    .p   (dSP_540_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_541 (
    .a   (dSP_541_a[7:0] ), //i
    .d   (dSP_541_d[7:0] ), //i
    .b   (dSP_541_b[7:0] ), //i
    .p   (dSP_541_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_542 (
    .a   (dSP_542_a[7:0] ), //i
    .d   (dSP_542_d[7:0] ), //i
    .b   (dSP_542_b[7:0] ), //i
    .p   (dSP_542_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_543 (
    .a   (dSP_543_a[7:0] ), //i
    .d   (dSP_543_d[7:0] ), //i
    .b   (dSP_543_b[7:0] ), //i
    .p   (dSP_543_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_544 (
    .a   (dSP_544_a[7:0] ), //i
    .d   (dSP_544_d[7:0] ), //i
    .b   (dSP_544_b[7:0] ), //i
    .p   (dSP_544_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_545 (
    .a   (dSP_545_a[7:0] ), //i
    .d   (dSP_545_d[7:0] ), //i
    .b   (dSP_545_b[7:0] ), //i
    .p   (dSP_545_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_546 (
    .a   (dSP_546_a[7:0] ), //i
    .d   (dSP_546_d[7:0] ), //i
    .b   (dSP_546_b[7:0] ), //i
    .p   (dSP_546_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_547 (
    .a   (dSP_547_a[7:0] ), //i
    .d   (dSP_547_d[7:0] ), //i
    .b   (dSP_547_b[7:0] ), //i
    .p   (dSP_547_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_548 (
    .a   (dSP_548_a[7:0] ), //i
    .d   (dSP_548_d[7:0] ), //i
    .b   (dSP_548_b[7:0] ), //i
    .p   (dSP_548_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_549 (
    .a   (dSP_549_a[7:0] ), //i
    .d   (dSP_549_d[7:0] ), //i
    .b   (dSP_549_b[7:0] ), //i
    .p   (dSP_549_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_550 (
    .a   (dSP_550_a[7:0] ), //i
    .d   (dSP_550_d[7:0] ), //i
    .b   (dSP_550_b[7:0] ), //i
    .p   (dSP_550_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_551 (
    .a   (dSP_551_a[7:0] ), //i
    .d   (dSP_551_d[7:0] ), //i
    .b   (dSP_551_b[7:0] ), //i
    .p   (dSP_551_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_552 (
    .a   (dSP_552_a[7:0] ), //i
    .d   (dSP_552_d[7:0] ), //i
    .b   (dSP_552_b[7:0] ), //i
    .p   (dSP_552_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_553 (
    .a   (dSP_553_a[7:0] ), //i
    .d   (dSP_553_d[7:0] ), //i
    .b   (dSP_553_b[7:0] ), //i
    .p   (dSP_553_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_554 (
    .a   (dSP_554_a[7:0] ), //i
    .d   (dSP_554_d[7:0] ), //i
    .b   (dSP_554_b[7:0] ), //i
    .p   (dSP_554_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_555 (
    .a   (dSP_555_a[7:0] ), //i
    .d   (dSP_555_d[7:0] ), //i
    .b   (dSP_555_b[7:0] ), //i
    .p   (dSP_555_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_556 (
    .a   (dSP_556_a[7:0] ), //i
    .d   (dSP_556_d[7:0] ), //i
    .b   (dSP_556_b[7:0] ), //i
    .p   (dSP_556_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_557 (
    .a   (dSP_557_a[7:0] ), //i
    .d   (dSP_557_d[7:0] ), //i
    .b   (dSP_557_b[7:0] ), //i
    .p   (dSP_557_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_558 (
    .a   (dSP_558_a[7:0] ), //i
    .d   (dSP_558_d[7:0] ), //i
    .b   (dSP_558_b[7:0] ), //i
    .p   (dSP_558_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_559 (
    .a   (dSP_559_a[7:0] ), //i
    .d   (dSP_559_d[7:0] ), //i
    .b   (dSP_559_b[7:0] ), //i
    .p   (dSP_559_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_560 (
    .a   (dSP_560_a[7:0] ), //i
    .d   (dSP_560_d[7:0] ), //i
    .b   (dSP_560_b[7:0] ), //i
    .p   (dSP_560_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_561 (
    .a   (dSP_561_a[7:0] ), //i
    .d   (dSP_561_d[7:0] ), //i
    .b   (dSP_561_b[7:0] ), //i
    .p   (dSP_561_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_562 (
    .a   (dSP_562_a[7:0] ), //i
    .d   (dSP_562_d[7:0] ), //i
    .b   (dSP_562_b[7:0] ), //i
    .p   (dSP_562_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_563 (
    .a   (dSP_563_a[7:0] ), //i
    .d   (dSP_563_d[7:0] ), //i
    .b   (dSP_563_b[7:0] ), //i
    .p   (dSP_563_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_564 (
    .a   (dSP_564_a[7:0] ), //i
    .d   (dSP_564_d[7:0] ), //i
    .b   (dSP_564_b[7:0] ), //i
    .p   (dSP_564_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_565 (
    .a   (dSP_565_a[7:0] ), //i
    .d   (dSP_565_d[7:0] ), //i
    .b   (dSP_565_b[7:0] ), //i
    .p   (dSP_565_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_566 (
    .a   (dSP_566_a[7:0] ), //i
    .d   (dSP_566_d[7:0] ), //i
    .b   (dSP_566_b[7:0] ), //i
    .p   (dSP_566_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_567 (
    .a   (dSP_567_a[7:0] ), //i
    .d   (dSP_567_d[7:0] ), //i
    .b   (dSP_567_b[7:0] ), //i
    .p   (dSP_567_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_568 (
    .a   (dSP_568_a[7:0] ), //i
    .d   (dSP_568_d[7:0] ), //i
    .b   (dSP_568_b[7:0] ), //i
    .p   (dSP_568_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_569 (
    .a   (dSP_569_a[7:0] ), //i
    .d   (dSP_569_d[7:0] ), //i
    .b   (dSP_569_b[7:0] ), //i
    .p   (dSP_569_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_570 (
    .a   (dSP_570_a[7:0] ), //i
    .d   (dSP_570_d[7:0] ), //i
    .b   (dSP_570_b[7:0] ), //i
    .p   (dSP_570_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_571 (
    .a   (dSP_571_a[7:0] ), //i
    .d   (dSP_571_d[7:0] ), //i
    .b   (dSP_571_b[7:0] ), //i
    .p   (dSP_571_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_572 (
    .a   (dSP_572_a[7:0] ), //i
    .d   (dSP_572_d[7:0] ), //i
    .b   (dSP_572_b[7:0] ), //i
    .p   (dSP_572_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_573 (
    .a   (dSP_573_a[7:0] ), //i
    .d   (dSP_573_d[7:0] ), //i
    .b   (dSP_573_b[7:0] ), //i
    .p   (dSP_573_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_574 (
    .a   (dSP_574_a[7:0] ), //i
    .d   (dSP_574_d[7:0] ), //i
    .b   (dSP_574_b[7:0] ), //i
    .p   (dSP_574_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_575 (
    .a   (dSP_575_a[7:0] ), //i
    .d   (dSP_575_d[7:0] ), //i
    .b   (dSP_575_b[7:0] ), //i
    .p   (dSP_575_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_576 (
    .a   (dSP_576_a[7:0] ), //i
    .d   (dSP_576_d[7:0] ), //i
    .b   (dSP_576_b[7:0] ), //i
    .p   (dSP_576_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_577 (
    .a   (dSP_577_a[7:0] ), //i
    .d   (dSP_577_d[7:0] ), //i
    .b   (dSP_577_b[7:0] ), //i
    .p   (dSP_577_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_578 (
    .a   (dSP_578_a[7:0] ), //i
    .d   (dSP_578_d[7:0] ), //i
    .b   (dSP_578_b[7:0] ), //i
    .p   (dSP_578_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_579 (
    .a   (dSP_579_a[7:0] ), //i
    .d   (dSP_579_d[7:0] ), //i
    .b   (dSP_579_b[7:0] ), //i
    .p   (dSP_579_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_580 (
    .a   (dSP_580_a[7:0] ), //i
    .d   (dSP_580_d[7:0] ), //i
    .b   (dSP_580_b[7:0] ), //i
    .p   (dSP_580_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_581 (
    .a   (dSP_581_a[7:0] ), //i
    .d   (dSP_581_d[7:0] ), //i
    .b   (dSP_581_b[7:0] ), //i
    .p   (dSP_581_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_582 (
    .a   (dSP_582_a[7:0] ), //i
    .d   (dSP_582_d[7:0] ), //i
    .b   (dSP_582_b[7:0] ), //i
    .p   (dSP_582_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_583 (
    .a   (dSP_583_a[7:0] ), //i
    .d   (dSP_583_d[7:0] ), //i
    .b   (dSP_583_b[7:0] ), //i
    .p   (dSP_583_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_584 (
    .a   (dSP_584_a[7:0] ), //i
    .d   (dSP_584_d[7:0] ), //i
    .b   (dSP_584_b[7:0] ), //i
    .p   (dSP_584_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_585 (
    .a   (dSP_585_a[7:0] ), //i
    .d   (dSP_585_d[7:0] ), //i
    .b   (dSP_585_b[7:0] ), //i
    .p   (dSP_585_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_586 (
    .a   (dSP_586_a[7:0] ), //i
    .d   (dSP_586_d[7:0] ), //i
    .b   (dSP_586_b[7:0] ), //i
    .p   (dSP_586_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_587 (
    .a   (dSP_587_a[7:0] ), //i
    .d   (dSP_587_d[7:0] ), //i
    .b   (dSP_587_b[7:0] ), //i
    .p   (dSP_587_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_588 (
    .a   (dSP_588_a[7:0] ), //i
    .d   (dSP_588_d[7:0] ), //i
    .b   (dSP_588_b[7:0] ), //i
    .p   (dSP_588_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_589 (
    .a   (dSP_589_a[7:0] ), //i
    .d   (dSP_589_d[7:0] ), //i
    .b   (dSP_589_b[7:0] ), //i
    .p   (dSP_589_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_590 (
    .a   (dSP_590_a[7:0] ), //i
    .d   (dSP_590_d[7:0] ), //i
    .b   (dSP_590_b[7:0] ), //i
    .p   (dSP_590_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_591 (
    .a   (dSP_591_a[7:0] ), //i
    .d   (dSP_591_d[7:0] ), //i
    .b   (dSP_591_b[7:0] ), //i
    .p   (dSP_591_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_592 (
    .a   (dSP_592_a[7:0] ), //i
    .d   (dSP_592_d[7:0] ), //i
    .b   (dSP_592_b[7:0] ), //i
    .p   (dSP_592_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_593 (
    .a   (dSP_593_a[7:0] ), //i
    .d   (dSP_593_d[7:0] ), //i
    .b   (dSP_593_b[7:0] ), //i
    .p   (dSP_593_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_594 (
    .a   (dSP_594_a[7:0] ), //i
    .d   (dSP_594_d[7:0] ), //i
    .b   (dSP_594_b[7:0] ), //i
    .p   (dSP_594_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_595 (
    .a   (dSP_595_a[7:0] ), //i
    .d   (dSP_595_d[7:0] ), //i
    .b   (dSP_595_b[7:0] ), //i
    .p   (dSP_595_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_596 (
    .a   (dSP_596_a[7:0] ), //i
    .d   (dSP_596_d[7:0] ), //i
    .b   (dSP_596_b[7:0] ), //i
    .p   (dSP_596_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_597 (
    .a   (dSP_597_a[7:0] ), //i
    .d   (dSP_597_d[7:0] ), //i
    .b   (dSP_597_b[7:0] ), //i
    .p   (dSP_597_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_598 (
    .a   (dSP_598_a[7:0] ), //i
    .d   (dSP_598_d[7:0] ), //i
    .b   (dSP_598_b[7:0] ), //i
    .p   (dSP_598_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_599 (
    .a   (dSP_599_a[7:0] ), //i
    .d   (dSP_599_d[7:0] ), //i
    .b   (dSP_599_b[7:0] ), //i
    .p   (dSP_599_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_600 (
    .a   (dSP_600_a[7:0] ), //i
    .d   (dSP_600_d[7:0] ), //i
    .b   (dSP_600_b[7:0] ), //i
    .p   (dSP_600_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_601 (
    .a   (dSP_601_a[7:0] ), //i
    .d   (dSP_601_d[7:0] ), //i
    .b   (dSP_601_b[7:0] ), //i
    .p   (dSP_601_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_602 (
    .a   (dSP_602_a[7:0] ), //i
    .d   (dSP_602_d[7:0] ), //i
    .b   (dSP_602_b[7:0] ), //i
    .p   (dSP_602_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_603 (
    .a   (dSP_603_a[7:0] ), //i
    .d   (dSP_603_d[7:0] ), //i
    .b   (dSP_603_b[7:0] ), //i
    .p   (dSP_603_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_604 (
    .a   (dSP_604_a[7:0] ), //i
    .d   (dSP_604_d[7:0] ), //i
    .b   (dSP_604_b[7:0] ), //i
    .p   (dSP_604_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_605 (
    .a   (dSP_605_a[7:0] ), //i
    .d   (dSP_605_d[7:0] ), //i
    .b   (dSP_605_b[7:0] ), //i
    .p   (dSP_605_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_606 (
    .a   (dSP_606_a[7:0] ), //i
    .d   (dSP_606_d[7:0] ), //i
    .b   (dSP_606_b[7:0] ), //i
    .p   (dSP_606_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_607 (
    .a   (dSP_607_a[7:0] ), //i
    .d   (dSP_607_d[7:0] ), //i
    .b   (dSP_607_b[7:0] ), //i
    .p   (dSP_607_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_608 (
    .a   (dSP_608_a[7:0] ), //i
    .d   (dSP_608_d[7:0] ), //i
    .b   (dSP_608_b[7:0] ), //i
    .p   (dSP_608_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_609 (
    .a   (dSP_609_a[7:0] ), //i
    .d   (dSP_609_d[7:0] ), //i
    .b   (dSP_609_b[7:0] ), //i
    .p   (dSP_609_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_610 (
    .a   (dSP_610_a[7:0] ), //i
    .d   (dSP_610_d[7:0] ), //i
    .b   (dSP_610_b[7:0] ), //i
    .p   (dSP_610_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_611 (
    .a   (dSP_611_a[7:0] ), //i
    .d   (dSP_611_d[7:0] ), //i
    .b   (dSP_611_b[7:0] ), //i
    .p   (dSP_611_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_612 (
    .a   (dSP_612_a[7:0] ), //i
    .d   (dSP_612_d[7:0] ), //i
    .b   (dSP_612_b[7:0] ), //i
    .p   (dSP_612_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_613 (
    .a   (dSP_613_a[7:0] ), //i
    .d   (dSP_613_d[7:0] ), //i
    .b   (dSP_613_b[7:0] ), //i
    .p   (dSP_613_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_614 (
    .a   (dSP_614_a[7:0] ), //i
    .d   (dSP_614_d[7:0] ), //i
    .b   (dSP_614_b[7:0] ), //i
    .p   (dSP_614_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_615 (
    .a   (dSP_615_a[7:0] ), //i
    .d   (dSP_615_d[7:0] ), //i
    .b   (dSP_615_b[7:0] ), //i
    .p   (dSP_615_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_616 (
    .a   (dSP_616_a[7:0] ), //i
    .d   (dSP_616_d[7:0] ), //i
    .b   (dSP_616_b[7:0] ), //i
    .p   (dSP_616_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_617 (
    .a   (dSP_617_a[7:0] ), //i
    .d   (dSP_617_d[7:0] ), //i
    .b   (dSP_617_b[7:0] ), //i
    .p   (dSP_617_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_618 (
    .a   (dSP_618_a[7:0] ), //i
    .d   (dSP_618_d[7:0] ), //i
    .b   (dSP_618_b[7:0] ), //i
    .p   (dSP_618_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_619 (
    .a   (dSP_619_a[7:0] ), //i
    .d   (dSP_619_d[7:0] ), //i
    .b   (dSP_619_b[7:0] ), //i
    .p   (dSP_619_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_620 (
    .a   (dSP_620_a[7:0] ), //i
    .d   (dSP_620_d[7:0] ), //i
    .b   (dSP_620_b[7:0] ), //i
    .p   (dSP_620_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_621 (
    .a   (dSP_621_a[7:0] ), //i
    .d   (dSP_621_d[7:0] ), //i
    .b   (dSP_621_b[7:0] ), //i
    .p   (dSP_621_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_622 (
    .a   (dSP_622_a[7:0] ), //i
    .d   (dSP_622_d[7:0] ), //i
    .b   (dSP_622_b[7:0] ), //i
    .p   (dSP_622_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_623 (
    .a   (dSP_623_a[7:0] ), //i
    .d   (dSP_623_d[7:0] ), //i
    .b   (dSP_623_b[7:0] ), //i
    .p   (dSP_623_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_624 (
    .a   (dSP_624_a[7:0] ), //i
    .d   (dSP_624_d[7:0] ), //i
    .b   (dSP_624_b[7:0] ), //i
    .p   (dSP_624_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_625 (
    .a   (dSP_625_a[7:0] ), //i
    .d   (dSP_625_d[7:0] ), //i
    .b   (dSP_625_b[7:0] ), //i
    .p   (dSP_625_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_626 (
    .a   (dSP_626_a[7:0] ), //i
    .d   (dSP_626_d[7:0] ), //i
    .b   (dSP_626_b[7:0] ), //i
    .p   (dSP_626_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_627 (
    .a   (dSP_627_a[7:0] ), //i
    .d   (dSP_627_d[7:0] ), //i
    .b   (dSP_627_b[7:0] ), //i
    .p   (dSP_627_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_628 (
    .a   (dSP_628_a[7:0] ), //i
    .d   (dSP_628_d[7:0] ), //i
    .b   (dSP_628_b[7:0] ), //i
    .p   (dSP_628_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_629 (
    .a   (dSP_629_a[7:0] ), //i
    .d   (dSP_629_d[7:0] ), //i
    .b   (dSP_629_b[7:0] ), //i
    .p   (dSP_629_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_630 (
    .a   (dSP_630_a[7:0] ), //i
    .d   (dSP_630_d[7:0] ), //i
    .b   (dSP_630_b[7:0] ), //i
    .p   (dSP_630_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_631 (
    .a   (dSP_631_a[7:0] ), //i
    .d   (dSP_631_d[7:0] ), //i
    .b   (dSP_631_b[7:0] ), //i
    .p   (dSP_631_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_632 (
    .a   (dSP_632_a[7:0] ), //i
    .d   (dSP_632_d[7:0] ), //i
    .b   (dSP_632_b[7:0] ), //i
    .p   (dSP_632_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_633 (
    .a   (dSP_633_a[7:0] ), //i
    .d   (dSP_633_d[7:0] ), //i
    .b   (dSP_633_b[7:0] ), //i
    .p   (dSP_633_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_634 (
    .a   (dSP_634_a[7:0] ), //i
    .d   (dSP_634_d[7:0] ), //i
    .b   (dSP_634_b[7:0] ), //i
    .p   (dSP_634_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_635 (
    .a   (dSP_635_a[7:0] ), //i
    .d   (dSP_635_d[7:0] ), //i
    .b   (dSP_635_b[7:0] ), //i
    .p   (dSP_635_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_636 (
    .a   (dSP_636_a[7:0] ), //i
    .d   (dSP_636_d[7:0] ), //i
    .b   (dSP_636_b[7:0] ), //i
    .p   (dSP_636_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_637 (
    .a   (dSP_637_a[7:0] ), //i
    .d   (dSP_637_d[7:0] ), //i
    .b   (dSP_637_b[7:0] ), //i
    .p   (dSP_637_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_638 (
    .a   (dSP_638_a[7:0] ), //i
    .d   (dSP_638_d[7:0] ), //i
    .b   (dSP_638_b[7:0] ), //i
    .p   (dSP_638_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_639 (
    .a   (dSP_639_a[7:0] ), //i
    .d   (dSP_639_d[7:0] ), //i
    .b   (dSP_639_b[7:0] ), //i
    .p   (dSP_639_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_640 (
    .a   (dSP_640_a[7:0] ), //i
    .d   (dSP_640_d[7:0] ), //i
    .b   (dSP_640_b[7:0] ), //i
    .p   (dSP_640_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_641 (
    .a   (dSP_641_a[7:0] ), //i
    .d   (dSP_641_d[7:0] ), //i
    .b   (dSP_641_b[7:0] ), //i
    .p   (dSP_641_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_642 (
    .a   (dSP_642_a[7:0] ), //i
    .d   (dSP_642_d[7:0] ), //i
    .b   (dSP_642_b[7:0] ), //i
    .p   (dSP_642_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_643 (
    .a   (dSP_643_a[7:0] ), //i
    .d   (dSP_643_d[7:0] ), //i
    .b   (dSP_643_b[7:0] ), //i
    .p   (dSP_643_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_644 (
    .a   (dSP_644_a[7:0] ), //i
    .d   (dSP_644_d[7:0] ), //i
    .b   (dSP_644_b[7:0] ), //i
    .p   (dSP_644_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_645 (
    .a   (dSP_645_a[7:0] ), //i
    .d   (dSP_645_d[7:0] ), //i
    .b   (dSP_645_b[7:0] ), //i
    .p   (dSP_645_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_646 (
    .a   (dSP_646_a[7:0] ), //i
    .d   (dSP_646_d[7:0] ), //i
    .b   (dSP_646_b[7:0] ), //i
    .p   (dSP_646_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_647 (
    .a   (dSP_647_a[7:0] ), //i
    .d   (dSP_647_d[7:0] ), //i
    .b   (dSP_647_b[7:0] ), //i
    .p   (dSP_647_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_648 (
    .a   (dSP_648_a[7:0] ), //i
    .d   (dSP_648_d[7:0] ), //i
    .b   (dSP_648_b[7:0] ), //i
    .p   (dSP_648_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_649 (
    .a   (dSP_649_a[7:0] ), //i
    .d   (dSP_649_d[7:0] ), //i
    .b   (dSP_649_b[7:0] ), //i
    .p   (dSP_649_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_650 (
    .a   (dSP_650_a[7:0] ), //i
    .d   (dSP_650_d[7:0] ), //i
    .b   (dSP_650_b[7:0] ), //i
    .p   (dSP_650_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_651 (
    .a   (dSP_651_a[7:0] ), //i
    .d   (dSP_651_d[7:0] ), //i
    .b   (dSP_651_b[7:0] ), //i
    .p   (dSP_651_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_652 (
    .a   (dSP_652_a[7:0] ), //i
    .d   (dSP_652_d[7:0] ), //i
    .b   (dSP_652_b[7:0] ), //i
    .p   (dSP_652_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_653 (
    .a   (dSP_653_a[7:0] ), //i
    .d   (dSP_653_d[7:0] ), //i
    .b   (dSP_653_b[7:0] ), //i
    .p   (dSP_653_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_654 (
    .a   (dSP_654_a[7:0] ), //i
    .d   (dSP_654_d[7:0] ), //i
    .b   (dSP_654_b[7:0] ), //i
    .p   (dSP_654_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_655 (
    .a   (dSP_655_a[7:0] ), //i
    .d   (dSP_655_d[7:0] ), //i
    .b   (dSP_655_b[7:0] ), //i
    .p   (dSP_655_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_656 (
    .a   (dSP_656_a[7:0] ), //i
    .d   (dSP_656_d[7:0] ), //i
    .b   (dSP_656_b[7:0] ), //i
    .p   (dSP_656_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_657 (
    .a   (dSP_657_a[7:0] ), //i
    .d   (dSP_657_d[7:0] ), //i
    .b   (dSP_657_b[7:0] ), //i
    .p   (dSP_657_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_658 (
    .a   (dSP_658_a[7:0] ), //i
    .d   (dSP_658_d[7:0] ), //i
    .b   (dSP_658_b[7:0] ), //i
    .p   (dSP_658_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_659 (
    .a   (dSP_659_a[7:0] ), //i
    .d   (dSP_659_d[7:0] ), //i
    .b   (dSP_659_b[7:0] ), //i
    .p   (dSP_659_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_660 (
    .a   (dSP_660_a[7:0] ), //i
    .d   (dSP_660_d[7:0] ), //i
    .b   (dSP_660_b[7:0] ), //i
    .p   (dSP_660_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_661 (
    .a   (dSP_661_a[7:0] ), //i
    .d   (dSP_661_d[7:0] ), //i
    .b   (dSP_661_b[7:0] ), //i
    .p   (dSP_661_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_662 (
    .a   (dSP_662_a[7:0] ), //i
    .d   (dSP_662_d[7:0] ), //i
    .b   (dSP_662_b[7:0] ), //i
    .p   (dSP_662_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_663 (
    .a   (dSP_663_a[7:0] ), //i
    .d   (dSP_663_d[7:0] ), //i
    .b   (dSP_663_b[7:0] ), //i
    .p   (dSP_663_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_664 (
    .a   (dSP_664_a[7:0] ), //i
    .d   (dSP_664_d[7:0] ), //i
    .b   (dSP_664_b[7:0] ), //i
    .p   (dSP_664_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_665 (
    .a   (dSP_665_a[7:0] ), //i
    .d   (dSP_665_d[7:0] ), //i
    .b   (dSP_665_b[7:0] ), //i
    .p   (dSP_665_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_666 (
    .a   (dSP_666_a[7:0] ), //i
    .d   (dSP_666_d[7:0] ), //i
    .b   (dSP_666_b[7:0] ), //i
    .p   (dSP_666_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_667 (
    .a   (dSP_667_a[7:0] ), //i
    .d   (dSP_667_d[7:0] ), //i
    .b   (dSP_667_b[7:0] ), //i
    .p   (dSP_667_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_668 (
    .a   (dSP_668_a[7:0] ), //i
    .d   (dSP_668_d[7:0] ), //i
    .b   (dSP_668_b[7:0] ), //i
    .p   (dSP_668_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_669 (
    .a   (dSP_669_a[7:0] ), //i
    .d   (dSP_669_d[7:0] ), //i
    .b   (dSP_669_b[7:0] ), //i
    .p   (dSP_669_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_670 (
    .a   (dSP_670_a[7:0] ), //i
    .d   (dSP_670_d[7:0] ), //i
    .b   (dSP_670_b[7:0] ), //i
    .p   (dSP_670_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_671 (
    .a   (dSP_671_a[7:0] ), //i
    .d   (dSP_671_d[7:0] ), //i
    .b   (dSP_671_b[7:0] ), //i
    .p   (dSP_671_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_672 (
    .a   (dSP_672_a[7:0] ), //i
    .d   (dSP_672_d[7:0] ), //i
    .b   (dSP_672_b[7:0] ), //i
    .p   (dSP_672_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_673 (
    .a   (dSP_673_a[7:0] ), //i
    .d   (dSP_673_d[7:0] ), //i
    .b   (dSP_673_b[7:0] ), //i
    .p   (dSP_673_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_674 (
    .a   (dSP_674_a[7:0] ), //i
    .d   (dSP_674_d[7:0] ), //i
    .b   (dSP_674_b[7:0] ), //i
    .p   (dSP_674_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_675 (
    .a   (dSP_675_a[7:0] ), //i
    .d   (dSP_675_d[7:0] ), //i
    .b   (dSP_675_b[7:0] ), //i
    .p   (dSP_675_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_676 (
    .a   (dSP_676_a[7:0] ), //i
    .d   (dSP_676_d[7:0] ), //i
    .b   (dSP_676_b[7:0] ), //i
    .p   (dSP_676_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_677 (
    .a   (dSP_677_a[7:0] ), //i
    .d   (dSP_677_d[7:0] ), //i
    .b   (dSP_677_b[7:0] ), //i
    .p   (dSP_677_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_678 (
    .a   (dSP_678_a[7:0] ), //i
    .d   (dSP_678_d[7:0] ), //i
    .b   (dSP_678_b[7:0] ), //i
    .p   (dSP_678_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_679 (
    .a   (dSP_679_a[7:0] ), //i
    .d   (dSP_679_d[7:0] ), //i
    .b   (dSP_679_b[7:0] ), //i
    .p   (dSP_679_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_680 (
    .a   (dSP_680_a[7:0] ), //i
    .d   (dSP_680_d[7:0] ), //i
    .b   (dSP_680_b[7:0] ), //i
    .p   (dSP_680_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_681 (
    .a   (dSP_681_a[7:0] ), //i
    .d   (dSP_681_d[7:0] ), //i
    .b   (dSP_681_b[7:0] ), //i
    .p   (dSP_681_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_682 (
    .a   (dSP_682_a[7:0] ), //i
    .d   (dSP_682_d[7:0] ), //i
    .b   (dSP_682_b[7:0] ), //i
    .p   (dSP_682_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_683 (
    .a   (dSP_683_a[7:0] ), //i
    .d   (dSP_683_d[7:0] ), //i
    .b   (dSP_683_b[7:0] ), //i
    .p   (dSP_683_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_684 (
    .a   (dSP_684_a[7:0] ), //i
    .d   (dSP_684_d[7:0] ), //i
    .b   (dSP_684_b[7:0] ), //i
    .p   (dSP_684_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_685 (
    .a   (dSP_685_a[7:0] ), //i
    .d   (dSP_685_d[7:0] ), //i
    .b   (dSP_685_b[7:0] ), //i
    .p   (dSP_685_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_686 (
    .a   (dSP_686_a[7:0] ), //i
    .d   (dSP_686_d[7:0] ), //i
    .b   (dSP_686_b[7:0] ), //i
    .p   (dSP_686_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_687 (
    .a   (dSP_687_a[7:0] ), //i
    .d   (dSP_687_d[7:0] ), //i
    .b   (dSP_687_b[7:0] ), //i
    .p   (dSP_687_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_688 (
    .a   (dSP_688_a[7:0] ), //i
    .d   (dSP_688_d[7:0] ), //i
    .b   (dSP_688_b[7:0] ), //i
    .p   (dSP_688_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_689 (
    .a   (dSP_689_a[7:0] ), //i
    .d   (dSP_689_d[7:0] ), //i
    .b   (dSP_689_b[7:0] ), //i
    .p   (dSP_689_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_690 (
    .a   (dSP_690_a[7:0] ), //i
    .d   (dSP_690_d[7:0] ), //i
    .b   (dSP_690_b[7:0] ), //i
    .p   (dSP_690_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_691 (
    .a   (dSP_691_a[7:0] ), //i
    .d   (dSP_691_d[7:0] ), //i
    .b   (dSP_691_b[7:0] ), //i
    .p   (dSP_691_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_692 (
    .a   (dSP_692_a[7:0] ), //i
    .d   (dSP_692_d[7:0] ), //i
    .b   (dSP_692_b[7:0] ), //i
    .p   (dSP_692_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_693 (
    .a   (dSP_693_a[7:0] ), //i
    .d   (dSP_693_d[7:0] ), //i
    .b   (dSP_693_b[7:0] ), //i
    .p   (dSP_693_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_694 (
    .a   (dSP_694_a[7:0] ), //i
    .d   (dSP_694_d[7:0] ), //i
    .b   (dSP_694_b[7:0] ), //i
    .p   (dSP_694_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_695 (
    .a   (dSP_695_a[7:0] ), //i
    .d   (dSP_695_d[7:0] ), //i
    .b   (dSP_695_b[7:0] ), //i
    .p   (dSP_695_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_696 (
    .a   (dSP_696_a[7:0] ), //i
    .d   (dSP_696_d[7:0] ), //i
    .b   (dSP_696_b[7:0] ), //i
    .p   (dSP_696_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_697 (
    .a   (dSP_697_a[7:0] ), //i
    .d   (dSP_697_d[7:0] ), //i
    .b   (dSP_697_b[7:0] ), //i
    .p   (dSP_697_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_698 (
    .a   (dSP_698_a[7:0] ), //i
    .d   (dSP_698_d[7:0] ), //i
    .b   (dSP_698_b[7:0] ), //i
    .p   (dSP_698_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_699 (
    .a   (dSP_699_a[7:0] ), //i
    .d   (dSP_699_d[7:0] ), //i
    .b   (dSP_699_b[7:0] ), //i
    .p   (dSP_699_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_700 (
    .a   (dSP_700_a[7:0] ), //i
    .d   (dSP_700_d[7:0] ), //i
    .b   (dSP_700_b[7:0] ), //i
    .p   (dSP_700_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_701 (
    .a   (dSP_701_a[7:0] ), //i
    .d   (dSP_701_d[7:0] ), //i
    .b   (dSP_701_b[7:0] ), //i
    .p   (dSP_701_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_702 (
    .a   (dSP_702_a[7:0] ), //i
    .d   (dSP_702_d[7:0] ), //i
    .b   (dSP_702_b[7:0] ), //i
    .p   (dSP_702_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_703 (
    .a   (dSP_703_a[7:0] ), //i
    .d   (dSP_703_d[7:0] ), //i
    .b   (dSP_703_b[7:0] ), //i
    .p   (dSP_703_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_704 (
    .a   (dSP_704_a[7:0] ), //i
    .d   (dSP_704_d[7:0] ), //i
    .b   (dSP_704_b[7:0] ), //i
    .p   (dSP_704_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_705 (
    .a   (dSP_705_a[7:0] ), //i
    .d   (dSP_705_d[7:0] ), //i
    .b   (dSP_705_b[7:0] ), //i
    .p   (dSP_705_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_706 (
    .a   (dSP_706_a[7:0] ), //i
    .d   (dSP_706_d[7:0] ), //i
    .b   (dSP_706_b[7:0] ), //i
    .p   (dSP_706_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_707 (
    .a   (dSP_707_a[7:0] ), //i
    .d   (dSP_707_d[7:0] ), //i
    .b   (dSP_707_b[7:0] ), //i
    .p   (dSP_707_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_708 (
    .a   (dSP_708_a[7:0] ), //i
    .d   (dSP_708_d[7:0] ), //i
    .b   (dSP_708_b[7:0] ), //i
    .p   (dSP_708_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_709 (
    .a   (dSP_709_a[7:0] ), //i
    .d   (dSP_709_d[7:0] ), //i
    .b   (dSP_709_b[7:0] ), //i
    .p   (dSP_709_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_710 (
    .a   (dSP_710_a[7:0] ), //i
    .d   (dSP_710_d[7:0] ), //i
    .b   (dSP_710_b[7:0] ), //i
    .p   (dSP_710_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_711 (
    .a   (dSP_711_a[7:0] ), //i
    .d   (dSP_711_d[7:0] ), //i
    .b   (dSP_711_b[7:0] ), //i
    .p   (dSP_711_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_712 (
    .a   (dSP_712_a[7:0] ), //i
    .d   (dSP_712_d[7:0] ), //i
    .b   (dSP_712_b[7:0] ), //i
    .p   (dSP_712_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_713 (
    .a   (dSP_713_a[7:0] ), //i
    .d   (dSP_713_d[7:0] ), //i
    .b   (dSP_713_b[7:0] ), //i
    .p   (dSP_713_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_714 (
    .a   (dSP_714_a[7:0] ), //i
    .d   (dSP_714_d[7:0] ), //i
    .b   (dSP_714_b[7:0] ), //i
    .p   (dSP_714_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_715 (
    .a   (dSP_715_a[7:0] ), //i
    .d   (dSP_715_d[7:0] ), //i
    .b   (dSP_715_b[7:0] ), //i
    .p   (dSP_715_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_716 (
    .a   (dSP_716_a[7:0] ), //i
    .d   (dSP_716_d[7:0] ), //i
    .b   (dSP_716_b[7:0] ), //i
    .p   (dSP_716_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_717 (
    .a   (dSP_717_a[7:0] ), //i
    .d   (dSP_717_d[7:0] ), //i
    .b   (dSP_717_b[7:0] ), //i
    .p   (dSP_717_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_718 (
    .a   (dSP_718_a[7:0] ), //i
    .d   (dSP_718_d[7:0] ), //i
    .b   (dSP_718_b[7:0] ), //i
    .p   (dSP_718_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_719 (
    .a   (dSP_719_a[7:0] ), //i
    .d   (dSP_719_d[7:0] ), //i
    .b   (dSP_719_b[7:0] ), //i
    .p   (dSP_719_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_720 (
    .a   (dSP_720_a[7:0] ), //i
    .d   (dSP_720_d[7:0] ), //i
    .b   (dSP_720_b[7:0] ), //i
    .p   (dSP_720_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_721 (
    .a   (dSP_721_a[7:0] ), //i
    .d   (dSP_721_d[7:0] ), //i
    .b   (dSP_721_b[7:0] ), //i
    .p   (dSP_721_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_722 (
    .a   (dSP_722_a[7:0] ), //i
    .d   (dSP_722_d[7:0] ), //i
    .b   (dSP_722_b[7:0] ), //i
    .p   (dSP_722_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_723 (
    .a   (dSP_723_a[7:0] ), //i
    .d   (dSP_723_d[7:0] ), //i
    .b   (dSP_723_b[7:0] ), //i
    .p   (dSP_723_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_724 (
    .a   (dSP_724_a[7:0] ), //i
    .d   (dSP_724_d[7:0] ), //i
    .b   (dSP_724_b[7:0] ), //i
    .p   (dSP_724_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_725 (
    .a   (dSP_725_a[7:0] ), //i
    .d   (dSP_725_d[7:0] ), //i
    .b   (dSP_725_b[7:0] ), //i
    .p   (dSP_725_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_726 (
    .a   (dSP_726_a[7:0] ), //i
    .d   (dSP_726_d[7:0] ), //i
    .b   (dSP_726_b[7:0] ), //i
    .p   (dSP_726_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_727 (
    .a   (dSP_727_a[7:0] ), //i
    .d   (dSP_727_d[7:0] ), //i
    .b   (dSP_727_b[7:0] ), //i
    .p   (dSP_727_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_728 (
    .a   (dSP_728_a[7:0] ), //i
    .d   (dSP_728_d[7:0] ), //i
    .b   (dSP_728_b[7:0] ), //i
    .p   (dSP_728_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_729 (
    .a   (dSP_729_a[7:0] ), //i
    .d   (dSP_729_d[7:0] ), //i
    .b   (dSP_729_b[7:0] ), //i
    .p   (dSP_729_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_730 (
    .a   (dSP_730_a[7:0] ), //i
    .d   (dSP_730_d[7:0] ), //i
    .b   (dSP_730_b[7:0] ), //i
    .p   (dSP_730_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_731 (
    .a   (dSP_731_a[7:0] ), //i
    .d   (dSP_731_d[7:0] ), //i
    .b   (dSP_731_b[7:0] ), //i
    .p   (dSP_731_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_732 (
    .a   (dSP_732_a[7:0] ), //i
    .d   (dSP_732_d[7:0] ), //i
    .b   (dSP_732_b[7:0] ), //i
    .p   (dSP_732_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_733 (
    .a   (dSP_733_a[7:0] ), //i
    .d   (dSP_733_d[7:0] ), //i
    .b   (dSP_733_b[7:0] ), //i
    .p   (dSP_733_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_734 (
    .a   (dSP_734_a[7:0] ), //i
    .d   (dSP_734_d[7:0] ), //i
    .b   (dSP_734_b[7:0] ), //i
    .p   (dSP_734_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_735 (
    .a   (dSP_735_a[7:0] ), //i
    .d   (dSP_735_d[7:0] ), //i
    .b   (dSP_735_b[7:0] ), //i
    .p   (dSP_735_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_736 (
    .a   (dSP_736_a[7:0] ), //i
    .d   (dSP_736_d[7:0] ), //i
    .b   (dSP_736_b[7:0] ), //i
    .p   (dSP_736_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_737 (
    .a   (dSP_737_a[7:0] ), //i
    .d   (dSP_737_d[7:0] ), //i
    .b   (dSP_737_b[7:0] ), //i
    .p   (dSP_737_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_738 (
    .a   (dSP_738_a[7:0] ), //i
    .d   (dSP_738_d[7:0] ), //i
    .b   (dSP_738_b[7:0] ), //i
    .p   (dSP_738_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_739 (
    .a   (dSP_739_a[7:0] ), //i
    .d   (dSP_739_d[7:0] ), //i
    .b   (dSP_739_b[7:0] ), //i
    .p   (dSP_739_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_740 (
    .a   (dSP_740_a[7:0] ), //i
    .d   (dSP_740_d[7:0] ), //i
    .b   (dSP_740_b[7:0] ), //i
    .p   (dSP_740_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_741 (
    .a   (dSP_741_a[7:0] ), //i
    .d   (dSP_741_d[7:0] ), //i
    .b   (dSP_741_b[7:0] ), //i
    .p   (dSP_741_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_742 (
    .a   (dSP_742_a[7:0] ), //i
    .d   (dSP_742_d[7:0] ), //i
    .b   (dSP_742_b[7:0] ), //i
    .p   (dSP_742_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_743 (
    .a   (dSP_743_a[7:0] ), //i
    .d   (dSP_743_d[7:0] ), //i
    .b   (dSP_743_b[7:0] ), //i
    .p   (dSP_743_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_744 (
    .a   (dSP_744_a[7:0] ), //i
    .d   (dSP_744_d[7:0] ), //i
    .b   (dSP_744_b[7:0] ), //i
    .p   (dSP_744_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_745 (
    .a   (dSP_745_a[7:0] ), //i
    .d   (dSP_745_d[7:0] ), //i
    .b   (dSP_745_b[7:0] ), //i
    .p   (dSP_745_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_746 (
    .a   (dSP_746_a[7:0] ), //i
    .d   (dSP_746_d[7:0] ), //i
    .b   (dSP_746_b[7:0] ), //i
    .p   (dSP_746_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_747 (
    .a   (dSP_747_a[7:0] ), //i
    .d   (dSP_747_d[7:0] ), //i
    .b   (dSP_747_b[7:0] ), //i
    .p   (dSP_747_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_748 (
    .a   (dSP_748_a[7:0] ), //i
    .d   (dSP_748_d[7:0] ), //i
    .b   (dSP_748_b[7:0] ), //i
    .p   (dSP_748_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_749 (
    .a   (dSP_749_a[7:0] ), //i
    .d   (dSP_749_d[7:0] ), //i
    .b   (dSP_749_b[7:0] ), //i
    .p   (dSP_749_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_750 (
    .a   (dSP_750_a[7:0] ), //i
    .d   (dSP_750_d[7:0] ), //i
    .b   (dSP_750_b[7:0] ), //i
    .p   (dSP_750_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_751 (
    .a   (dSP_751_a[7:0] ), //i
    .d   (dSP_751_d[7:0] ), //i
    .b   (dSP_751_b[7:0] ), //i
    .p   (dSP_751_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_752 (
    .a   (dSP_752_a[7:0] ), //i
    .d   (dSP_752_d[7:0] ), //i
    .b   (dSP_752_b[7:0] ), //i
    .p   (dSP_752_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_753 (
    .a   (dSP_753_a[7:0] ), //i
    .d   (dSP_753_d[7:0] ), //i
    .b   (dSP_753_b[7:0] ), //i
    .p   (dSP_753_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_754 (
    .a   (dSP_754_a[7:0] ), //i
    .d   (dSP_754_d[7:0] ), //i
    .b   (dSP_754_b[7:0] ), //i
    .p   (dSP_754_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_755 (
    .a   (dSP_755_a[7:0] ), //i
    .d   (dSP_755_d[7:0] ), //i
    .b   (dSP_755_b[7:0] ), //i
    .p   (dSP_755_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_756 (
    .a   (dSP_756_a[7:0] ), //i
    .d   (dSP_756_d[7:0] ), //i
    .b   (dSP_756_b[7:0] ), //i
    .p   (dSP_756_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_757 (
    .a   (dSP_757_a[7:0] ), //i
    .d   (dSP_757_d[7:0] ), //i
    .b   (dSP_757_b[7:0] ), //i
    .p   (dSP_757_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_758 (
    .a   (dSP_758_a[7:0] ), //i
    .d   (dSP_758_d[7:0] ), //i
    .b   (dSP_758_b[7:0] ), //i
    .p   (dSP_758_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_759 (
    .a   (dSP_759_a[7:0] ), //i
    .d   (dSP_759_d[7:0] ), //i
    .b   (dSP_759_b[7:0] ), //i
    .p   (dSP_759_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_760 (
    .a   (dSP_760_a[7:0] ), //i
    .d   (dSP_760_d[7:0] ), //i
    .b   (dSP_760_b[7:0] ), //i
    .p   (dSP_760_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_761 (
    .a   (dSP_761_a[7:0] ), //i
    .d   (dSP_761_d[7:0] ), //i
    .b   (dSP_761_b[7:0] ), //i
    .p   (dSP_761_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_762 (
    .a   (dSP_762_a[7:0] ), //i
    .d   (dSP_762_d[7:0] ), //i
    .b   (dSP_762_b[7:0] ), //i
    .p   (dSP_762_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_763 (
    .a   (dSP_763_a[7:0] ), //i
    .d   (dSP_763_d[7:0] ), //i
    .b   (dSP_763_b[7:0] ), //i
    .p   (dSP_763_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_764 (
    .a   (dSP_764_a[7:0] ), //i
    .d   (dSP_764_d[7:0] ), //i
    .b   (dSP_764_b[7:0] ), //i
    .p   (dSP_764_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_765 (
    .a   (dSP_765_a[7:0] ), //i
    .d   (dSP_765_d[7:0] ), //i
    .b   (dSP_765_b[7:0] ), //i
    .p   (dSP_765_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_766 (
    .a   (dSP_766_a[7:0] ), //i
    .d   (dSP_766_d[7:0] ), //i
    .b   (dSP_766_b[7:0] ), //i
    .p   (dSP_766_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_767 (
    .a   (dSP_767_a[7:0] ), //i
    .d   (dSP_767_d[7:0] ), //i
    .b   (dSP_767_b[7:0] ), //i
    .p   (dSP_767_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_768 (
    .a   (dSP_768_a[7:0] ), //i
    .d   (dSP_768_d[7:0] ), //i
    .b   (dSP_768_b[7:0] ), //i
    .p   (dSP_768_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_769 (
    .a   (dSP_769_a[7:0] ), //i
    .d   (dSP_769_d[7:0] ), //i
    .b   (dSP_769_b[7:0] ), //i
    .p   (dSP_769_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_770 (
    .a   (dSP_770_a[7:0] ), //i
    .d   (dSP_770_d[7:0] ), //i
    .b   (dSP_770_b[7:0] ), //i
    .p   (dSP_770_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_771 (
    .a   (dSP_771_a[7:0] ), //i
    .d   (dSP_771_d[7:0] ), //i
    .b   (dSP_771_b[7:0] ), //i
    .p   (dSP_771_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_772 (
    .a   (dSP_772_a[7:0] ), //i
    .d   (dSP_772_d[7:0] ), //i
    .b   (dSP_772_b[7:0] ), //i
    .p   (dSP_772_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_773 (
    .a   (dSP_773_a[7:0] ), //i
    .d   (dSP_773_d[7:0] ), //i
    .b   (dSP_773_b[7:0] ), //i
    .p   (dSP_773_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_774 (
    .a   (dSP_774_a[7:0] ), //i
    .d   (dSP_774_d[7:0] ), //i
    .b   (dSP_774_b[7:0] ), //i
    .p   (dSP_774_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_775 (
    .a   (dSP_775_a[7:0] ), //i
    .d   (dSP_775_d[7:0] ), //i
    .b   (dSP_775_b[7:0] ), //i
    .p   (dSP_775_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_776 (
    .a   (dSP_776_a[7:0] ), //i
    .d   (dSP_776_d[7:0] ), //i
    .b   (dSP_776_b[7:0] ), //i
    .p   (dSP_776_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_777 (
    .a   (dSP_777_a[7:0] ), //i
    .d   (dSP_777_d[7:0] ), //i
    .b   (dSP_777_b[7:0] ), //i
    .p   (dSP_777_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_778 (
    .a   (dSP_778_a[7:0] ), //i
    .d   (dSP_778_d[7:0] ), //i
    .b   (dSP_778_b[7:0] ), //i
    .p   (dSP_778_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_779 (
    .a   (dSP_779_a[7:0] ), //i
    .d   (dSP_779_d[7:0] ), //i
    .b   (dSP_779_b[7:0] ), //i
    .p   (dSP_779_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_780 (
    .a   (dSP_780_a[7:0] ), //i
    .d   (dSP_780_d[7:0] ), //i
    .b   (dSP_780_b[7:0] ), //i
    .p   (dSP_780_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_781 (
    .a   (dSP_781_a[7:0] ), //i
    .d   (dSP_781_d[7:0] ), //i
    .b   (dSP_781_b[7:0] ), //i
    .p   (dSP_781_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_782 (
    .a   (dSP_782_a[7:0] ), //i
    .d   (dSP_782_d[7:0] ), //i
    .b   (dSP_782_b[7:0] ), //i
    .p   (dSP_782_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_783 (
    .a   (dSP_783_a[7:0] ), //i
    .d   (dSP_783_d[7:0] ), //i
    .b   (dSP_783_b[7:0] ), //i
    .p   (dSP_783_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_784 (
    .a   (dSP_784_a[7:0] ), //i
    .d   (dSP_784_d[7:0] ), //i
    .b   (dSP_784_b[7:0] ), //i
    .p   (dSP_784_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_785 (
    .a   (dSP_785_a[7:0] ), //i
    .d   (dSP_785_d[7:0] ), //i
    .b   (dSP_785_b[7:0] ), //i
    .p   (dSP_785_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_786 (
    .a   (dSP_786_a[7:0] ), //i
    .d   (dSP_786_d[7:0] ), //i
    .b   (dSP_786_b[7:0] ), //i
    .p   (dSP_786_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_787 (
    .a   (dSP_787_a[7:0] ), //i
    .d   (dSP_787_d[7:0] ), //i
    .b   (dSP_787_b[7:0] ), //i
    .p   (dSP_787_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_788 (
    .a   (dSP_788_a[7:0] ), //i
    .d   (dSP_788_d[7:0] ), //i
    .b   (dSP_788_b[7:0] ), //i
    .p   (dSP_788_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_789 (
    .a   (dSP_789_a[7:0] ), //i
    .d   (dSP_789_d[7:0] ), //i
    .b   (dSP_789_b[7:0] ), //i
    .p   (dSP_789_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_790 (
    .a   (dSP_790_a[7:0] ), //i
    .d   (dSP_790_d[7:0] ), //i
    .b   (dSP_790_b[7:0] ), //i
    .p   (dSP_790_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_791 (
    .a   (dSP_791_a[7:0] ), //i
    .d   (dSP_791_d[7:0] ), //i
    .b   (dSP_791_b[7:0] ), //i
    .p   (dSP_791_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_792 (
    .a   (dSP_792_a[7:0] ), //i
    .d   (dSP_792_d[7:0] ), //i
    .b   (dSP_792_b[7:0] ), //i
    .p   (dSP_792_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_793 (
    .a   (dSP_793_a[7:0] ), //i
    .d   (dSP_793_d[7:0] ), //i
    .b   (dSP_793_b[7:0] ), //i
    .p   (dSP_793_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_794 (
    .a   (dSP_794_a[7:0] ), //i
    .d   (dSP_794_d[7:0] ), //i
    .b   (dSP_794_b[7:0] ), //i
    .p   (dSP_794_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_795 (
    .a   (dSP_795_a[7:0] ), //i
    .d   (dSP_795_d[7:0] ), //i
    .b   (dSP_795_b[7:0] ), //i
    .p   (dSP_795_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_796 (
    .a   (dSP_796_a[7:0] ), //i
    .d   (dSP_796_d[7:0] ), //i
    .b   (dSP_796_b[7:0] ), //i
    .p   (dSP_796_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_797 (
    .a   (dSP_797_a[7:0] ), //i
    .d   (dSP_797_d[7:0] ), //i
    .b   (dSP_797_b[7:0] ), //i
    .p   (dSP_797_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_798 (
    .a   (dSP_798_a[7:0] ), //i
    .d   (dSP_798_d[7:0] ), //i
    .b   (dSP_798_b[7:0] ), //i
    .p   (dSP_798_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_799 (
    .a   (dSP_799_a[7:0] ), //i
    .d   (dSP_799_d[7:0] ), //i
    .b   (dSP_799_b[7:0] ), //i
    .p   (dSP_799_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_800 (
    .a   (dSP_800_a[7:0] ), //i
    .d   (dSP_800_d[7:0] ), //i
    .b   (dSP_800_b[7:0] ), //i
    .p   (dSP_800_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_801 (
    .a   (dSP_801_a[7:0] ), //i
    .d   (dSP_801_d[7:0] ), //i
    .b   (dSP_801_b[7:0] ), //i
    .p   (dSP_801_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_802 (
    .a   (dSP_802_a[7:0] ), //i
    .d   (dSP_802_d[7:0] ), //i
    .b   (dSP_802_b[7:0] ), //i
    .p   (dSP_802_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_803 (
    .a   (dSP_803_a[7:0] ), //i
    .d   (dSP_803_d[7:0] ), //i
    .b   (dSP_803_b[7:0] ), //i
    .p   (dSP_803_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_804 (
    .a   (dSP_804_a[7:0] ), //i
    .d   (dSP_804_d[7:0] ), //i
    .b   (dSP_804_b[7:0] ), //i
    .p   (dSP_804_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_805 (
    .a   (dSP_805_a[7:0] ), //i
    .d   (dSP_805_d[7:0] ), //i
    .b   (dSP_805_b[7:0] ), //i
    .p   (dSP_805_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_806 (
    .a   (dSP_806_a[7:0] ), //i
    .d   (dSP_806_d[7:0] ), //i
    .b   (dSP_806_b[7:0] ), //i
    .p   (dSP_806_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_807 (
    .a   (dSP_807_a[7:0] ), //i
    .d   (dSP_807_d[7:0] ), //i
    .b   (dSP_807_b[7:0] ), //i
    .p   (dSP_807_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_808 (
    .a   (dSP_808_a[7:0] ), //i
    .d   (dSP_808_d[7:0] ), //i
    .b   (dSP_808_b[7:0] ), //i
    .p   (dSP_808_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_809 (
    .a   (dSP_809_a[7:0] ), //i
    .d   (dSP_809_d[7:0] ), //i
    .b   (dSP_809_b[7:0] ), //i
    .p   (dSP_809_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_810 (
    .a   (dSP_810_a[7:0] ), //i
    .d   (dSP_810_d[7:0] ), //i
    .b   (dSP_810_b[7:0] ), //i
    .p   (dSP_810_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_811 (
    .a   (dSP_811_a[7:0] ), //i
    .d   (dSP_811_d[7:0] ), //i
    .b   (dSP_811_b[7:0] ), //i
    .p   (dSP_811_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_812 (
    .a   (dSP_812_a[7:0] ), //i
    .d   (dSP_812_d[7:0] ), //i
    .b   (dSP_812_b[7:0] ), //i
    .p   (dSP_812_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_813 (
    .a   (dSP_813_a[7:0] ), //i
    .d   (dSP_813_d[7:0] ), //i
    .b   (dSP_813_b[7:0] ), //i
    .p   (dSP_813_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_814 (
    .a   (dSP_814_a[7:0] ), //i
    .d   (dSP_814_d[7:0] ), //i
    .b   (dSP_814_b[7:0] ), //i
    .p   (dSP_814_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_815 (
    .a   (dSP_815_a[7:0] ), //i
    .d   (dSP_815_d[7:0] ), //i
    .b   (dSP_815_b[7:0] ), //i
    .p   (dSP_815_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_816 (
    .a   (dSP_816_a[7:0] ), //i
    .d   (dSP_816_d[7:0] ), //i
    .b   (dSP_816_b[7:0] ), //i
    .p   (dSP_816_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_817 (
    .a   (dSP_817_a[7:0] ), //i
    .d   (dSP_817_d[7:0] ), //i
    .b   (dSP_817_b[7:0] ), //i
    .p   (dSP_817_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_818 (
    .a   (dSP_818_a[7:0] ), //i
    .d   (dSP_818_d[7:0] ), //i
    .b   (dSP_818_b[7:0] ), //i
    .p   (dSP_818_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_819 (
    .a   (dSP_819_a[7:0] ), //i
    .d   (dSP_819_d[7:0] ), //i
    .b   (dSP_819_b[7:0] ), //i
    .p   (dSP_819_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_820 (
    .a   (dSP_820_a[7:0] ), //i
    .d   (dSP_820_d[7:0] ), //i
    .b   (dSP_820_b[7:0] ), //i
    .p   (dSP_820_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_821 (
    .a   (dSP_821_a[7:0] ), //i
    .d   (dSP_821_d[7:0] ), //i
    .b   (dSP_821_b[7:0] ), //i
    .p   (dSP_821_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_822 (
    .a   (dSP_822_a[7:0] ), //i
    .d   (dSP_822_d[7:0] ), //i
    .b   (dSP_822_b[7:0] ), //i
    .p   (dSP_822_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_823 (
    .a   (dSP_823_a[7:0] ), //i
    .d   (dSP_823_d[7:0] ), //i
    .b   (dSP_823_b[7:0] ), //i
    .p   (dSP_823_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_824 (
    .a   (dSP_824_a[7:0] ), //i
    .d   (dSP_824_d[7:0] ), //i
    .b   (dSP_824_b[7:0] ), //i
    .p   (dSP_824_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_825 (
    .a   (dSP_825_a[7:0] ), //i
    .d   (dSP_825_d[7:0] ), //i
    .b   (dSP_825_b[7:0] ), //i
    .p   (dSP_825_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_826 (
    .a   (dSP_826_a[7:0] ), //i
    .d   (dSP_826_d[7:0] ), //i
    .b   (dSP_826_b[7:0] ), //i
    .p   (dSP_826_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_827 (
    .a   (dSP_827_a[7:0] ), //i
    .d   (dSP_827_d[7:0] ), //i
    .b   (dSP_827_b[7:0] ), //i
    .p   (dSP_827_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_828 (
    .a   (dSP_828_a[7:0] ), //i
    .d   (dSP_828_d[7:0] ), //i
    .b   (dSP_828_b[7:0] ), //i
    .p   (dSP_828_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_829 (
    .a   (dSP_829_a[7:0] ), //i
    .d   (dSP_829_d[7:0] ), //i
    .b   (dSP_829_b[7:0] ), //i
    .p   (dSP_829_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_830 (
    .a   (dSP_830_a[7:0] ), //i
    .d   (dSP_830_d[7:0] ), //i
    .b   (dSP_830_b[7:0] ), //i
    .p   (dSP_830_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_831 (
    .a   (dSP_831_a[7:0] ), //i
    .d   (dSP_831_d[7:0] ), //i
    .b   (dSP_831_b[7:0] ), //i
    .p   (dSP_831_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_832 (
    .a   (dSP_832_a[7:0] ), //i
    .d   (dSP_832_d[7:0] ), //i
    .b   (dSP_832_b[7:0] ), //i
    .p   (dSP_832_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_833 (
    .a   (dSP_833_a[7:0] ), //i
    .d   (dSP_833_d[7:0] ), //i
    .b   (dSP_833_b[7:0] ), //i
    .p   (dSP_833_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_834 (
    .a   (dSP_834_a[7:0] ), //i
    .d   (dSP_834_d[7:0] ), //i
    .b   (dSP_834_b[7:0] ), //i
    .p   (dSP_834_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_835 (
    .a   (dSP_835_a[7:0] ), //i
    .d   (dSP_835_d[7:0] ), //i
    .b   (dSP_835_b[7:0] ), //i
    .p   (dSP_835_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_836 (
    .a   (dSP_836_a[7:0] ), //i
    .d   (dSP_836_d[7:0] ), //i
    .b   (dSP_836_b[7:0] ), //i
    .p   (dSP_836_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_837 (
    .a   (dSP_837_a[7:0] ), //i
    .d   (dSP_837_d[7:0] ), //i
    .b   (dSP_837_b[7:0] ), //i
    .p   (dSP_837_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_838 (
    .a   (dSP_838_a[7:0] ), //i
    .d   (dSP_838_d[7:0] ), //i
    .b   (dSP_838_b[7:0] ), //i
    .p   (dSP_838_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_839 (
    .a   (dSP_839_a[7:0] ), //i
    .d   (dSP_839_d[7:0] ), //i
    .b   (dSP_839_b[7:0] ), //i
    .p   (dSP_839_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_840 (
    .a   (dSP_840_a[7:0] ), //i
    .d   (dSP_840_d[7:0] ), //i
    .b   (dSP_840_b[7:0] ), //i
    .p   (dSP_840_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_841 (
    .a   (dSP_841_a[7:0] ), //i
    .d   (dSP_841_d[7:0] ), //i
    .b   (dSP_841_b[7:0] ), //i
    .p   (dSP_841_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_842 (
    .a   (dSP_842_a[7:0] ), //i
    .d   (dSP_842_d[7:0] ), //i
    .b   (dSP_842_b[7:0] ), //i
    .p   (dSP_842_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_843 (
    .a   (dSP_843_a[7:0] ), //i
    .d   (dSP_843_d[7:0] ), //i
    .b   (dSP_843_b[7:0] ), //i
    .p   (dSP_843_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_844 (
    .a   (dSP_844_a[7:0] ), //i
    .d   (dSP_844_d[7:0] ), //i
    .b   (dSP_844_b[7:0] ), //i
    .p   (dSP_844_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_845 (
    .a   (dSP_845_a[7:0] ), //i
    .d   (dSP_845_d[7:0] ), //i
    .b   (dSP_845_b[7:0] ), //i
    .p   (dSP_845_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_846 (
    .a   (dSP_846_a[7:0] ), //i
    .d   (dSP_846_d[7:0] ), //i
    .b   (dSP_846_b[7:0] ), //i
    .p   (dSP_846_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_847 (
    .a   (dSP_847_a[7:0] ), //i
    .d   (dSP_847_d[7:0] ), //i
    .b   (dSP_847_b[7:0] ), //i
    .p   (dSP_847_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_848 (
    .a   (dSP_848_a[7:0] ), //i
    .d   (dSP_848_d[7:0] ), //i
    .b   (dSP_848_b[7:0] ), //i
    .p   (dSP_848_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_849 (
    .a   (dSP_849_a[7:0] ), //i
    .d   (dSP_849_d[7:0] ), //i
    .b   (dSP_849_b[7:0] ), //i
    .p   (dSP_849_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_850 (
    .a   (dSP_850_a[7:0] ), //i
    .d   (dSP_850_d[7:0] ), //i
    .b   (dSP_850_b[7:0] ), //i
    .p   (dSP_850_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_851 (
    .a   (dSP_851_a[7:0] ), //i
    .d   (dSP_851_d[7:0] ), //i
    .b   (dSP_851_b[7:0] ), //i
    .p   (dSP_851_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_852 (
    .a   (dSP_852_a[7:0] ), //i
    .d   (dSP_852_d[7:0] ), //i
    .b   (dSP_852_b[7:0] ), //i
    .p   (dSP_852_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_853 (
    .a   (dSP_853_a[7:0] ), //i
    .d   (dSP_853_d[7:0] ), //i
    .b   (dSP_853_b[7:0] ), //i
    .p   (dSP_853_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_854 (
    .a   (dSP_854_a[7:0] ), //i
    .d   (dSP_854_d[7:0] ), //i
    .b   (dSP_854_b[7:0] ), //i
    .p   (dSP_854_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_855 (
    .a   (dSP_855_a[7:0] ), //i
    .d   (dSP_855_d[7:0] ), //i
    .b   (dSP_855_b[7:0] ), //i
    .p   (dSP_855_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_856 (
    .a   (dSP_856_a[7:0] ), //i
    .d   (dSP_856_d[7:0] ), //i
    .b   (dSP_856_b[7:0] ), //i
    .p   (dSP_856_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_857 (
    .a   (dSP_857_a[7:0] ), //i
    .d   (dSP_857_d[7:0] ), //i
    .b   (dSP_857_b[7:0] ), //i
    .p   (dSP_857_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_858 (
    .a   (dSP_858_a[7:0] ), //i
    .d   (dSP_858_d[7:0] ), //i
    .b   (dSP_858_b[7:0] ), //i
    .p   (dSP_858_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_859 (
    .a   (dSP_859_a[7:0] ), //i
    .d   (dSP_859_d[7:0] ), //i
    .b   (dSP_859_b[7:0] ), //i
    .p   (dSP_859_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_860 (
    .a   (dSP_860_a[7:0] ), //i
    .d   (dSP_860_d[7:0] ), //i
    .b   (dSP_860_b[7:0] ), //i
    .p   (dSP_860_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_861 (
    .a   (dSP_861_a[7:0] ), //i
    .d   (dSP_861_d[7:0] ), //i
    .b   (dSP_861_b[7:0] ), //i
    .p   (dSP_861_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_862 (
    .a   (dSP_862_a[7:0] ), //i
    .d   (dSP_862_d[7:0] ), //i
    .b   (dSP_862_b[7:0] ), //i
    .p   (dSP_862_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_863 (
    .a   (dSP_863_a[7:0] ), //i
    .d   (dSP_863_d[7:0] ), //i
    .b   (dSP_863_b[7:0] ), //i
    .p   (dSP_863_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_864 (
    .a   (dSP_864_a[7:0] ), //i
    .d   (dSP_864_d[7:0] ), //i
    .b   (dSP_864_b[7:0] ), //i
    .p   (dSP_864_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_865 (
    .a   (dSP_865_a[7:0] ), //i
    .d   (dSP_865_d[7:0] ), //i
    .b   (dSP_865_b[7:0] ), //i
    .p   (dSP_865_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_866 (
    .a   (dSP_866_a[7:0] ), //i
    .d   (dSP_866_d[7:0] ), //i
    .b   (dSP_866_b[7:0] ), //i
    .p   (dSP_866_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_867 (
    .a   (dSP_867_a[7:0] ), //i
    .d   (dSP_867_d[7:0] ), //i
    .b   (dSP_867_b[7:0] ), //i
    .p   (dSP_867_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_868 (
    .a   (dSP_868_a[7:0] ), //i
    .d   (dSP_868_d[7:0] ), //i
    .b   (dSP_868_b[7:0] ), //i
    .p   (dSP_868_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_869 (
    .a   (dSP_869_a[7:0] ), //i
    .d   (dSP_869_d[7:0] ), //i
    .b   (dSP_869_b[7:0] ), //i
    .p   (dSP_869_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_870 (
    .a   (dSP_870_a[7:0] ), //i
    .d   (dSP_870_d[7:0] ), //i
    .b   (dSP_870_b[7:0] ), //i
    .p   (dSP_870_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_871 (
    .a   (dSP_871_a[7:0] ), //i
    .d   (dSP_871_d[7:0] ), //i
    .b   (dSP_871_b[7:0] ), //i
    .p   (dSP_871_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_872 (
    .a   (dSP_872_a[7:0] ), //i
    .d   (dSP_872_d[7:0] ), //i
    .b   (dSP_872_b[7:0] ), //i
    .p   (dSP_872_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_873 (
    .a   (dSP_873_a[7:0] ), //i
    .d   (dSP_873_d[7:0] ), //i
    .b   (dSP_873_b[7:0] ), //i
    .p   (dSP_873_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_874 (
    .a   (dSP_874_a[7:0] ), //i
    .d   (dSP_874_d[7:0] ), //i
    .b   (dSP_874_b[7:0] ), //i
    .p   (dSP_874_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_875 (
    .a   (dSP_875_a[7:0] ), //i
    .d   (dSP_875_d[7:0] ), //i
    .b   (dSP_875_b[7:0] ), //i
    .p   (dSP_875_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_876 (
    .a   (dSP_876_a[7:0] ), //i
    .d   (dSP_876_d[7:0] ), //i
    .b   (dSP_876_b[7:0] ), //i
    .p   (dSP_876_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_877 (
    .a   (dSP_877_a[7:0] ), //i
    .d   (dSP_877_d[7:0] ), //i
    .b   (dSP_877_b[7:0] ), //i
    .p   (dSP_877_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_878 (
    .a   (dSP_878_a[7:0] ), //i
    .d   (dSP_878_d[7:0] ), //i
    .b   (dSP_878_b[7:0] ), //i
    .p   (dSP_878_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_879 (
    .a   (dSP_879_a[7:0] ), //i
    .d   (dSP_879_d[7:0] ), //i
    .b   (dSP_879_b[7:0] ), //i
    .p   (dSP_879_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_880 (
    .a   (dSP_880_a[7:0] ), //i
    .d   (dSP_880_d[7:0] ), //i
    .b   (dSP_880_b[7:0] ), //i
    .p   (dSP_880_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_881 (
    .a   (dSP_881_a[7:0] ), //i
    .d   (dSP_881_d[7:0] ), //i
    .b   (dSP_881_b[7:0] ), //i
    .p   (dSP_881_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_882 (
    .a   (dSP_882_a[7:0] ), //i
    .d   (dSP_882_d[7:0] ), //i
    .b   (dSP_882_b[7:0] ), //i
    .p   (dSP_882_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_883 (
    .a   (dSP_883_a[7:0] ), //i
    .d   (dSP_883_d[7:0] ), //i
    .b   (dSP_883_b[7:0] ), //i
    .p   (dSP_883_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_884 (
    .a   (dSP_884_a[7:0] ), //i
    .d   (dSP_884_d[7:0] ), //i
    .b   (dSP_884_b[7:0] ), //i
    .p   (dSP_884_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_885 (
    .a   (dSP_885_a[7:0] ), //i
    .d   (dSP_885_d[7:0] ), //i
    .b   (dSP_885_b[7:0] ), //i
    .p   (dSP_885_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_886 (
    .a   (dSP_886_a[7:0] ), //i
    .d   (dSP_886_d[7:0] ), //i
    .b   (dSP_886_b[7:0] ), //i
    .p   (dSP_886_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_887 (
    .a   (dSP_887_a[7:0] ), //i
    .d   (dSP_887_d[7:0] ), //i
    .b   (dSP_887_b[7:0] ), //i
    .p   (dSP_887_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_888 (
    .a   (dSP_888_a[7:0] ), //i
    .d   (dSP_888_d[7:0] ), //i
    .b   (dSP_888_b[7:0] ), //i
    .p   (dSP_888_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_889 (
    .a   (dSP_889_a[7:0] ), //i
    .d   (dSP_889_d[7:0] ), //i
    .b   (dSP_889_b[7:0] ), //i
    .p   (dSP_889_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_890 (
    .a   (dSP_890_a[7:0] ), //i
    .d   (dSP_890_d[7:0] ), //i
    .b   (dSP_890_b[7:0] ), //i
    .p   (dSP_890_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_891 (
    .a   (dSP_891_a[7:0] ), //i
    .d   (dSP_891_d[7:0] ), //i
    .b   (dSP_891_b[7:0] ), //i
    .p   (dSP_891_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_892 (
    .a   (dSP_892_a[7:0] ), //i
    .d   (dSP_892_d[7:0] ), //i
    .b   (dSP_892_b[7:0] ), //i
    .p   (dSP_892_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_893 (
    .a   (dSP_893_a[7:0] ), //i
    .d   (dSP_893_d[7:0] ), //i
    .b   (dSP_893_b[7:0] ), //i
    .p   (dSP_893_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_894 (
    .a   (dSP_894_a[7:0] ), //i
    .d   (dSP_894_d[7:0] ), //i
    .b   (dSP_894_b[7:0] ), //i
    .p   (dSP_894_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_895 (
    .a   (dSP_895_a[7:0] ), //i
    .d   (dSP_895_d[7:0] ), //i
    .b   (dSP_895_b[7:0] ), //i
    .p   (dSP_895_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_896 (
    .a   (dSP_896_a[7:0] ), //i
    .d   (dSP_896_d[7:0] ), //i
    .b   (dSP_896_b[7:0] ), //i
    .p   (dSP_896_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_897 (
    .a   (dSP_897_a[7:0] ), //i
    .d   (dSP_897_d[7:0] ), //i
    .b   (dSP_897_b[7:0] ), //i
    .p   (dSP_897_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_898 (
    .a   (dSP_898_a[7:0] ), //i
    .d   (dSP_898_d[7:0] ), //i
    .b   (dSP_898_b[7:0] ), //i
    .p   (dSP_898_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_899 (
    .a   (dSP_899_a[7:0] ), //i
    .d   (dSP_899_d[7:0] ), //i
    .b   (dSP_899_b[7:0] ), //i
    .p   (dSP_899_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_900 (
    .a   (dSP_900_a[7:0] ), //i
    .d   (dSP_900_d[7:0] ), //i
    .b   (dSP_900_b[7:0] ), //i
    .p   (dSP_900_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_901 (
    .a   (dSP_901_a[7:0] ), //i
    .d   (dSP_901_d[7:0] ), //i
    .b   (dSP_901_b[7:0] ), //i
    .p   (dSP_901_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_902 (
    .a   (dSP_902_a[7:0] ), //i
    .d   (dSP_902_d[7:0] ), //i
    .b   (dSP_902_b[7:0] ), //i
    .p   (dSP_902_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_903 (
    .a   (dSP_903_a[7:0] ), //i
    .d   (dSP_903_d[7:0] ), //i
    .b   (dSP_903_b[7:0] ), //i
    .p   (dSP_903_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_904 (
    .a   (dSP_904_a[7:0] ), //i
    .d   (dSP_904_d[7:0] ), //i
    .b   (dSP_904_b[7:0] ), //i
    .p   (dSP_904_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_905 (
    .a   (dSP_905_a[7:0] ), //i
    .d   (dSP_905_d[7:0] ), //i
    .b   (dSP_905_b[7:0] ), //i
    .p   (dSP_905_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_906 (
    .a   (dSP_906_a[7:0] ), //i
    .d   (dSP_906_d[7:0] ), //i
    .b   (dSP_906_b[7:0] ), //i
    .p   (dSP_906_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_907 (
    .a   (dSP_907_a[7:0] ), //i
    .d   (dSP_907_d[7:0] ), //i
    .b   (dSP_907_b[7:0] ), //i
    .p   (dSP_907_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_908 (
    .a   (dSP_908_a[7:0] ), //i
    .d   (dSP_908_d[7:0] ), //i
    .b   (dSP_908_b[7:0] ), //i
    .p   (dSP_908_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_909 (
    .a   (dSP_909_a[7:0] ), //i
    .d   (dSP_909_d[7:0] ), //i
    .b   (dSP_909_b[7:0] ), //i
    .p   (dSP_909_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_910 (
    .a   (dSP_910_a[7:0] ), //i
    .d   (dSP_910_d[7:0] ), //i
    .b   (dSP_910_b[7:0] ), //i
    .p   (dSP_910_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_911 (
    .a   (dSP_911_a[7:0] ), //i
    .d   (dSP_911_d[7:0] ), //i
    .b   (dSP_911_b[7:0] ), //i
    .p   (dSP_911_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_912 (
    .a   (dSP_912_a[7:0] ), //i
    .d   (dSP_912_d[7:0] ), //i
    .b   (dSP_912_b[7:0] ), //i
    .p   (dSP_912_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_913 (
    .a   (dSP_913_a[7:0] ), //i
    .d   (dSP_913_d[7:0] ), //i
    .b   (dSP_913_b[7:0] ), //i
    .p   (dSP_913_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_914 (
    .a   (dSP_914_a[7:0] ), //i
    .d   (dSP_914_d[7:0] ), //i
    .b   (dSP_914_b[7:0] ), //i
    .p   (dSP_914_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_915 (
    .a   (dSP_915_a[7:0] ), //i
    .d   (dSP_915_d[7:0] ), //i
    .b   (dSP_915_b[7:0] ), //i
    .p   (dSP_915_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_916 (
    .a   (dSP_916_a[7:0] ), //i
    .d   (dSP_916_d[7:0] ), //i
    .b   (dSP_916_b[7:0] ), //i
    .p   (dSP_916_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_917 (
    .a   (dSP_917_a[7:0] ), //i
    .d   (dSP_917_d[7:0] ), //i
    .b   (dSP_917_b[7:0] ), //i
    .p   (dSP_917_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_918 (
    .a   (dSP_918_a[7:0] ), //i
    .d   (dSP_918_d[7:0] ), //i
    .b   (dSP_918_b[7:0] ), //i
    .p   (dSP_918_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_919 (
    .a   (dSP_919_a[7:0] ), //i
    .d   (dSP_919_d[7:0] ), //i
    .b   (dSP_919_b[7:0] ), //i
    .p   (dSP_919_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_920 (
    .a   (dSP_920_a[7:0] ), //i
    .d   (dSP_920_d[7:0] ), //i
    .b   (dSP_920_b[7:0] ), //i
    .p   (dSP_920_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_921 (
    .a   (dSP_921_a[7:0] ), //i
    .d   (dSP_921_d[7:0] ), //i
    .b   (dSP_921_b[7:0] ), //i
    .p   (dSP_921_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_922 (
    .a   (dSP_922_a[7:0] ), //i
    .d   (dSP_922_d[7:0] ), //i
    .b   (dSP_922_b[7:0] ), //i
    .p   (dSP_922_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_923 (
    .a   (dSP_923_a[7:0] ), //i
    .d   (dSP_923_d[7:0] ), //i
    .b   (dSP_923_b[7:0] ), //i
    .p   (dSP_923_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_924 (
    .a   (dSP_924_a[7:0] ), //i
    .d   (dSP_924_d[7:0] ), //i
    .b   (dSP_924_b[7:0] ), //i
    .p   (dSP_924_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_925 (
    .a   (dSP_925_a[7:0] ), //i
    .d   (dSP_925_d[7:0] ), //i
    .b   (dSP_925_b[7:0] ), //i
    .p   (dSP_925_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_926 (
    .a   (dSP_926_a[7:0] ), //i
    .d   (dSP_926_d[7:0] ), //i
    .b   (dSP_926_b[7:0] ), //i
    .p   (dSP_926_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_927 (
    .a   (dSP_927_a[7:0] ), //i
    .d   (dSP_927_d[7:0] ), //i
    .b   (dSP_927_b[7:0] ), //i
    .p   (dSP_927_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_928 (
    .a   (dSP_928_a[7:0] ), //i
    .d   (dSP_928_d[7:0] ), //i
    .b   (dSP_928_b[7:0] ), //i
    .p   (dSP_928_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_929 (
    .a   (dSP_929_a[7:0] ), //i
    .d   (dSP_929_d[7:0] ), //i
    .b   (dSP_929_b[7:0] ), //i
    .p   (dSP_929_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_930 (
    .a   (dSP_930_a[7:0] ), //i
    .d   (dSP_930_d[7:0] ), //i
    .b   (dSP_930_b[7:0] ), //i
    .p   (dSP_930_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_931 (
    .a   (dSP_931_a[7:0] ), //i
    .d   (dSP_931_d[7:0] ), //i
    .b   (dSP_931_b[7:0] ), //i
    .p   (dSP_931_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_932 (
    .a   (dSP_932_a[7:0] ), //i
    .d   (dSP_932_d[7:0] ), //i
    .b   (dSP_932_b[7:0] ), //i
    .p   (dSP_932_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_933 (
    .a   (dSP_933_a[7:0] ), //i
    .d   (dSP_933_d[7:0] ), //i
    .b   (dSP_933_b[7:0] ), //i
    .p   (dSP_933_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_934 (
    .a   (dSP_934_a[7:0] ), //i
    .d   (dSP_934_d[7:0] ), //i
    .b   (dSP_934_b[7:0] ), //i
    .p   (dSP_934_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_935 (
    .a   (dSP_935_a[7:0] ), //i
    .d   (dSP_935_d[7:0] ), //i
    .b   (dSP_935_b[7:0] ), //i
    .p   (dSP_935_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_936 (
    .a   (dSP_936_a[7:0] ), //i
    .d   (dSP_936_d[7:0] ), //i
    .b   (dSP_936_b[7:0] ), //i
    .p   (dSP_936_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_937 (
    .a   (dSP_937_a[7:0] ), //i
    .d   (dSP_937_d[7:0] ), //i
    .b   (dSP_937_b[7:0] ), //i
    .p   (dSP_937_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_938 (
    .a   (dSP_938_a[7:0] ), //i
    .d   (dSP_938_d[7:0] ), //i
    .b   (dSP_938_b[7:0] ), //i
    .p   (dSP_938_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_939 (
    .a   (dSP_939_a[7:0] ), //i
    .d   (dSP_939_d[7:0] ), //i
    .b   (dSP_939_b[7:0] ), //i
    .p   (dSP_939_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_940 (
    .a   (dSP_940_a[7:0] ), //i
    .d   (dSP_940_d[7:0] ), //i
    .b   (dSP_940_b[7:0] ), //i
    .p   (dSP_940_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_941 (
    .a   (dSP_941_a[7:0] ), //i
    .d   (dSP_941_d[7:0] ), //i
    .b   (dSP_941_b[7:0] ), //i
    .p   (dSP_941_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_942 (
    .a   (dSP_942_a[7:0] ), //i
    .d   (dSP_942_d[7:0] ), //i
    .b   (dSP_942_b[7:0] ), //i
    .p   (dSP_942_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_943 (
    .a   (dSP_943_a[7:0] ), //i
    .d   (dSP_943_d[7:0] ), //i
    .b   (dSP_943_b[7:0] ), //i
    .p   (dSP_943_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_944 (
    .a   (dSP_944_a[7:0] ), //i
    .d   (dSP_944_d[7:0] ), //i
    .b   (dSP_944_b[7:0] ), //i
    .p   (dSP_944_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_945 (
    .a   (dSP_945_a[7:0] ), //i
    .d   (dSP_945_d[7:0] ), //i
    .b   (dSP_945_b[7:0] ), //i
    .p   (dSP_945_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_946 (
    .a   (dSP_946_a[7:0] ), //i
    .d   (dSP_946_d[7:0] ), //i
    .b   (dSP_946_b[7:0] ), //i
    .p   (dSP_946_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_947 (
    .a   (dSP_947_a[7:0] ), //i
    .d   (dSP_947_d[7:0] ), //i
    .b   (dSP_947_b[7:0] ), //i
    .p   (dSP_947_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_948 (
    .a   (dSP_948_a[7:0] ), //i
    .d   (dSP_948_d[7:0] ), //i
    .b   (dSP_948_b[7:0] ), //i
    .p   (dSP_948_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_949 (
    .a   (dSP_949_a[7:0] ), //i
    .d   (dSP_949_d[7:0] ), //i
    .b   (dSP_949_b[7:0] ), //i
    .p   (dSP_949_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_950 (
    .a   (dSP_950_a[7:0] ), //i
    .d   (dSP_950_d[7:0] ), //i
    .b   (dSP_950_b[7:0] ), //i
    .p   (dSP_950_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_951 (
    .a   (dSP_951_a[7:0] ), //i
    .d   (dSP_951_d[7:0] ), //i
    .b   (dSP_951_b[7:0] ), //i
    .p   (dSP_951_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_952 (
    .a   (dSP_952_a[7:0] ), //i
    .d   (dSP_952_d[7:0] ), //i
    .b   (dSP_952_b[7:0] ), //i
    .p   (dSP_952_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_953 (
    .a   (dSP_953_a[7:0] ), //i
    .d   (dSP_953_d[7:0] ), //i
    .b   (dSP_953_b[7:0] ), //i
    .p   (dSP_953_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_954 (
    .a   (dSP_954_a[7:0] ), //i
    .d   (dSP_954_d[7:0] ), //i
    .b   (dSP_954_b[7:0] ), //i
    .p   (dSP_954_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_955 (
    .a   (dSP_955_a[7:0] ), //i
    .d   (dSP_955_d[7:0] ), //i
    .b   (dSP_955_b[7:0] ), //i
    .p   (dSP_955_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_956 (
    .a   (dSP_956_a[7:0] ), //i
    .d   (dSP_956_d[7:0] ), //i
    .b   (dSP_956_b[7:0] ), //i
    .p   (dSP_956_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_957 (
    .a   (dSP_957_a[7:0] ), //i
    .d   (dSP_957_d[7:0] ), //i
    .b   (dSP_957_b[7:0] ), //i
    .p   (dSP_957_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_958 (
    .a   (dSP_958_a[7:0] ), //i
    .d   (dSP_958_d[7:0] ), //i
    .b   (dSP_958_b[7:0] ), //i
    .p   (dSP_958_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_959 (
    .a   (dSP_959_a[7:0] ), //i
    .d   (dSP_959_d[7:0] ), //i
    .b   (dSP_959_b[7:0] ), //i
    .p   (dSP_959_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_960 (
    .a   (dSP_960_a[7:0] ), //i
    .d   (dSP_960_d[7:0] ), //i
    .b   (dSP_960_b[7:0] ), //i
    .p   (dSP_960_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_961 (
    .a   (dSP_961_a[7:0] ), //i
    .d   (dSP_961_d[7:0] ), //i
    .b   (dSP_961_b[7:0] ), //i
    .p   (dSP_961_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_962 (
    .a   (dSP_962_a[7:0] ), //i
    .d   (dSP_962_d[7:0] ), //i
    .b   (dSP_962_b[7:0] ), //i
    .p   (dSP_962_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_963 (
    .a   (dSP_963_a[7:0] ), //i
    .d   (dSP_963_d[7:0] ), //i
    .b   (dSP_963_b[7:0] ), //i
    .p   (dSP_963_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_964 (
    .a   (dSP_964_a[7:0] ), //i
    .d   (dSP_964_d[7:0] ), //i
    .b   (dSP_964_b[7:0] ), //i
    .p   (dSP_964_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_965 (
    .a   (dSP_965_a[7:0] ), //i
    .d   (dSP_965_d[7:0] ), //i
    .b   (dSP_965_b[7:0] ), //i
    .p   (dSP_965_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_966 (
    .a   (dSP_966_a[7:0] ), //i
    .d   (dSP_966_d[7:0] ), //i
    .b   (dSP_966_b[7:0] ), //i
    .p   (dSP_966_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_967 (
    .a   (dSP_967_a[7:0] ), //i
    .d   (dSP_967_d[7:0] ), //i
    .b   (dSP_967_b[7:0] ), //i
    .p   (dSP_967_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_968 (
    .a   (dSP_968_a[7:0] ), //i
    .d   (dSP_968_d[7:0] ), //i
    .b   (dSP_968_b[7:0] ), //i
    .p   (dSP_968_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_969 (
    .a   (dSP_969_a[7:0] ), //i
    .d   (dSP_969_d[7:0] ), //i
    .b   (dSP_969_b[7:0] ), //i
    .p   (dSP_969_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_970 (
    .a   (dSP_970_a[7:0] ), //i
    .d   (dSP_970_d[7:0] ), //i
    .b   (dSP_970_b[7:0] ), //i
    .p   (dSP_970_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_971 (
    .a   (dSP_971_a[7:0] ), //i
    .d   (dSP_971_d[7:0] ), //i
    .b   (dSP_971_b[7:0] ), //i
    .p   (dSP_971_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_972 (
    .a   (dSP_972_a[7:0] ), //i
    .d   (dSP_972_d[7:0] ), //i
    .b   (dSP_972_b[7:0] ), //i
    .p   (dSP_972_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_973 (
    .a   (dSP_973_a[7:0] ), //i
    .d   (dSP_973_d[7:0] ), //i
    .b   (dSP_973_b[7:0] ), //i
    .p   (dSP_973_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_974 (
    .a   (dSP_974_a[7:0] ), //i
    .d   (dSP_974_d[7:0] ), //i
    .b   (dSP_974_b[7:0] ), //i
    .p   (dSP_974_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_975 (
    .a   (dSP_975_a[7:0] ), //i
    .d   (dSP_975_d[7:0] ), //i
    .b   (dSP_975_b[7:0] ), //i
    .p   (dSP_975_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_976 (
    .a   (dSP_976_a[7:0] ), //i
    .d   (dSP_976_d[7:0] ), //i
    .b   (dSP_976_b[7:0] ), //i
    .p   (dSP_976_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_977 (
    .a   (dSP_977_a[7:0] ), //i
    .d   (dSP_977_d[7:0] ), //i
    .b   (dSP_977_b[7:0] ), //i
    .p   (dSP_977_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_978 (
    .a   (dSP_978_a[7:0] ), //i
    .d   (dSP_978_d[7:0] ), //i
    .b   (dSP_978_b[7:0] ), //i
    .p   (dSP_978_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_979 (
    .a   (dSP_979_a[7:0] ), //i
    .d   (dSP_979_d[7:0] ), //i
    .b   (dSP_979_b[7:0] ), //i
    .p   (dSP_979_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_980 (
    .a   (dSP_980_a[7:0] ), //i
    .d   (dSP_980_d[7:0] ), //i
    .b   (dSP_980_b[7:0] ), //i
    .p   (dSP_980_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_981 (
    .a   (dSP_981_a[7:0] ), //i
    .d   (dSP_981_d[7:0] ), //i
    .b   (dSP_981_b[7:0] ), //i
    .p   (dSP_981_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_982 (
    .a   (dSP_982_a[7:0] ), //i
    .d   (dSP_982_d[7:0] ), //i
    .b   (dSP_982_b[7:0] ), //i
    .p   (dSP_982_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_983 (
    .a   (dSP_983_a[7:0] ), //i
    .d   (dSP_983_d[7:0] ), //i
    .b   (dSP_983_b[7:0] ), //i
    .p   (dSP_983_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_984 (
    .a   (dSP_984_a[7:0] ), //i
    .d   (dSP_984_d[7:0] ), //i
    .b   (dSP_984_b[7:0] ), //i
    .p   (dSP_984_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_985 (
    .a   (dSP_985_a[7:0] ), //i
    .d   (dSP_985_d[7:0] ), //i
    .b   (dSP_985_b[7:0] ), //i
    .p   (dSP_985_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_986 (
    .a   (dSP_986_a[7:0] ), //i
    .d   (dSP_986_d[7:0] ), //i
    .b   (dSP_986_b[7:0] ), //i
    .p   (dSP_986_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_987 (
    .a   (dSP_987_a[7:0] ), //i
    .d   (dSP_987_d[7:0] ), //i
    .b   (dSP_987_b[7:0] ), //i
    .p   (dSP_987_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_988 (
    .a   (dSP_988_a[7:0] ), //i
    .d   (dSP_988_d[7:0] ), //i
    .b   (dSP_988_b[7:0] ), //i
    .p   (dSP_988_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_989 (
    .a   (dSP_989_a[7:0] ), //i
    .d   (dSP_989_d[7:0] ), //i
    .b   (dSP_989_b[7:0] ), //i
    .p   (dSP_989_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_990 (
    .a   (dSP_990_a[7:0] ), //i
    .d   (dSP_990_d[7:0] ), //i
    .b   (dSP_990_b[7:0] ), //i
    .p   (dSP_990_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_991 (
    .a   (dSP_991_a[7:0] ), //i
    .d   (dSP_991_d[7:0] ), //i
    .b   (dSP_991_b[7:0] ), //i
    .p   (dSP_991_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_992 (
    .a   (dSP_992_a[7:0] ), //i
    .d   (dSP_992_d[7:0] ), //i
    .b   (dSP_992_b[7:0] ), //i
    .p   (dSP_992_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_993 (
    .a   (dSP_993_a[7:0] ), //i
    .d   (dSP_993_d[7:0] ), //i
    .b   (dSP_993_b[7:0] ), //i
    .p   (dSP_993_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_994 (
    .a   (dSP_994_a[7:0] ), //i
    .d   (dSP_994_d[7:0] ), //i
    .b   (dSP_994_b[7:0] ), //i
    .p   (dSP_994_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_995 (
    .a   (dSP_995_a[7:0] ), //i
    .d   (dSP_995_d[7:0] ), //i
    .b   (dSP_995_b[7:0] ), //i
    .p   (dSP_995_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_996 (
    .a   (dSP_996_a[7:0] ), //i
    .d   (dSP_996_d[7:0] ), //i
    .b   (dSP_996_b[7:0] ), //i
    .p   (dSP_996_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_997 (
    .a   (dSP_997_a[7:0] ), //i
    .d   (dSP_997_d[7:0] ), //i
    .b   (dSP_997_b[7:0] ), //i
    .p   (dSP_997_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_998 (
    .a   (dSP_998_a[7:0] ), //i
    .d   (dSP_998_d[7:0] ), //i
    .b   (dSP_998_b[7:0] ), //i
    .p   (dSP_998_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_999 (
    .a   (dSP_999_a[7:0] ), //i
    .d   (dSP_999_d[7:0] ), //i
    .b   (dSP_999_b[7:0] ), //i
    .p   (dSP_999_p[31:0]), //o
    .CLK (clk            )  //i
  );
  DSP dSP_1000 (
    .a   (dSP_1000_a[7:0] ), //i
    .d   (dSP_1000_d[7:0] ), //i
    .b   (dSP_1000_b[7:0] ), //i
    .p   (dSP_1000_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1001 (
    .a   (dSP_1001_a[7:0] ), //i
    .d   (dSP_1001_d[7:0] ), //i
    .b   (dSP_1001_b[7:0] ), //i
    .p   (dSP_1001_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1002 (
    .a   (dSP_1002_a[7:0] ), //i
    .d   (dSP_1002_d[7:0] ), //i
    .b   (dSP_1002_b[7:0] ), //i
    .p   (dSP_1002_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1003 (
    .a   (dSP_1003_a[7:0] ), //i
    .d   (dSP_1003_d[7:0] ), //i
    .b   (dSP_1003_b[7:0] ), //i
    .p   (dSP_1003_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1004 (
    .a   (dSP_1004_a[7:0] ), //i
    .d   (dSP_1004_d[7:0] ), //i
    .b   (dSP_1004_b[7:0] ), //i
    .p   (dSP_1004_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1005 (
    .a   (dSP_1005_a[7:0] ), //i
    .d   (dSP_1005_d[7:0] ), //i
    .b   (dSP_1005_b[7:0] ), //i
    .p   (dSP_1005_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1006 (
    .a   (dSP_1006_a[7:0] ), //i
    .d   (dSP_1006_d[7:0] ), //i
    .b   (dSP_1006_b[7:0] ), //i
    .p   (dSP_1006_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1007 (
    .a   (dSP_1007_a[7:0] ), //i
    .d   (dSP_1007_d[7:0] ), //i
    .b   (dSP_1007_b[7:0] ), //i
    .p   (dSP_1007_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1008 (
    .a   (dSP_1008_a[7:0] ), //i
    .d   (dSP_1008_d[7:0] ), //i
    .b   (dSP_1008_b[7:0] ), //i
    .p   (dSP_1008_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1009 (
    .a   (dSP_1009_a[7:0] ), //i
    .d   (dSP_1009_d[7:0] ), //i
    .b   (dSP_1009_b[7:0] ), //i
    .p   (dSP_1009_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1010 (
    .a   (dSP_1010_a[7:0] ), //i
    .d   (dSP_1010_d[7:0] ), //i
    .b   (dSP_1010_b[7:0] ), //i
    .p   (dSP_1010_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1011 (
    .a   (dSP_1011_a[7:0] ), //i
    .d   (dSP_1011_d[7:0] ), //i
    .b   (dSP_1011_b[7:0] ), //i
    .p   (dSP_1011_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1012 (
    .a   (dSP_1012_a[7:0] ), //i
    .d   (dSP_1012_d[7:0] ), //i
    .b   (dSP_1012_b[7:0] ), //i
    .p   (dSP_1012_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1013 (
    .a   (dSP_1013_a[7:0] ), //i
    .d   (dSP_1013_d[7:0] ), //i
    .b   (dSP_1013_b[7:0] ), //i
    .p   (dSP_1013_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1014 (
    .a   (dSP_1014_a[7:0] ), //i
    .d   (dSP_1014_d[7:0] ), //i
    .b   (dSP_1014_b[7:0] ), //i
    .p   (dSP_1014_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1015 (
    .a   (dSP_1015_a[7:0] ), //i
    .d   (dSP_1015_d[7:0] ), //i
    .b   (dSP_1015_b[7:0] ), //i
    .p   (dSP_1015_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1016 (
    .a   (dSP_1016_a[7:0] ), //i
    .d   (dSP_1016_d[7:0] ), //i
    .b   (dSP_1016_b[7:0] ), //i
    .p   (dSP_1016_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1017 (
    .a   (dSP_1017_a[7:0] ), //i
    .d   (dSP_1017_d[7:0] ), //i
    .b   (dSP_1017_b[7:0] ), //i
    .p   (dSP_1017_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1018 (
    .a   (dSP_1018_a[7:0] ), //i
    .d   (dSP_1018_d[7:0] ), //i
    .b   (dSP_1018_b[7:0] ), //i
    .p   (dSP_1018_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1019 (
    .a   (dSP_1019_a[7:0] ), //i
    .d   (dSP_1019_d[7:0] ), //i
    .b   (dSP_1019_b[7:0] ), //i
    .p   (dSP_1019_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1020 (
    .a   (dSP_1020_a[7:0] ), //i
    .d   (dSP_1020_d[7:0] ), //i
    .b   (dSP_1020_b[7:0] ), //i
    .p   (dSP_1020_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1021 (
    .a   (dSP_1021_a[7:0] ), //i
    .d   (dSP_1021_d[7:0] ), //i
    .b   (dSP_1021_b[7:0] ), //i
    .p   (dSP_1021_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1022 (
    .a   (dSP_1022_a[7:0] ), //i
    .d   (dSP_1022_d[7:0] ), //i
    .b   (dSP_1022_b[7:0] ), //i
    .p   (dSP_1022_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1023 (
    .a   (dSP_1023_a[7:0] ), //i
    .d   (dSP_1023_d[7:0] ), //i
    .b   (dSP_1023_b[7:0] ), //i
    .p   (dSP_1023_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1024 (
    .a   (dSP_1024_a[7:0] ), //i
    .d   (dSP_1024_d[7:0] ), //i
    .b   (dSP_1024_b[7:0] ), //i
    .p   (dSP_1024_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1025 (
    .a   (dSP_1025_a[7:0] ), //i
    .d   (dSP_1025_d[7:0] ), //i
    .b   (dSP_1025_b[7:0] ), //i
    .p   (dSP_1025_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1026 (
    .a   (dSP_1026_a[7:0] ), //i
    .d   (dSP_1026_d[7:0] ), //i
    .b   (dSP_1026_b[7:0] ), //i
    .p   (dSP_1026_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1027 (
    .a   (dSP_1027_a[7:0] ), //i
    .d   (dSP_1027_d[7:0] ), //i
    .b   (dSP_1027_b[7:0] ), //i
    .p   (dSP_1027_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1028 (
    .a   (dSP_1028_a[7:0] ), //i
    .d   (dSP_1028_d[7:0] ), //i
    .b   (dSP_1028_b[7:0] ), //i
    .p   (dSP_1028_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1029 (
    .a   (dSP_1029_a[7:0] ), //i
    .d   (dSP_1029_d[7:0] ), //i
    .b   (dSP_1029_b[7:0] ), //i
    .p   (dSP_1029_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1030 (
    .a   (dSP_1030_a[7:0] ), //i
    .d   (dSP_1030_d[7:0] ), //i
    .b   (dSP_1030_b[7:0] ), //i
    .p   (dSP_1030_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1031 (
    .a   (dSP_1031_a[7:0] ), //i
    .d   (dSP_1031_d[7:0] ), //i
    .b   (dSP_1031_b[7:0] ), //i
    .p   (dSP_1031_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1032 (
    .a   (dSP_1032_a[7:0] ), //i
    .d   (dSP_1032_d[7:0] ), //i
    .b   (dSP_1032_b[7:0] ), //i
    .p   (dSP_1032_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1033 (
    .a   (dSP_1033_a[7:0] ), //i
    .d   (dSP_1033_d[7:0] ), //i
    .b   (dSP_1033_b[7:0] ), //i
    .p   (dSP_1033_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1034 (
    .a   (dSP_1034_a[7:0] ), //i
    .d   (dSP_1034_d[7:0] ), //i
    .b   (dSP_1034_b[7:0] ), //i
    .p   (dSP_1034_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1035 (
    .a   (dSP_1035_a[7:0] ), //i
    .d   (dSP_1035_d[7:0] ), //i
    .b   (dSP_1035_b[7:0] ), //i
    .p   (dSP_1035_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1036 (
    .a   (dSP_1036_a[7:0] ), //i
    .d   (dSP_1036_d[7:0] ), //i
    .b   (dSP_1036_b[7:0] ), //i
    .p   (dSP_1036_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1037 (
    .a   (dSP_1037_a[7:0] ), //i
    .d   (dSP_1037_d[7:0] ), //i
    .b   (dSP_1037_b[7:0] ), //i
    .p   (dSP_1037_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1038 (
    .a   (dSP_1038_a[7:0] ), //i
    .d   (dSP_1038_d[7:0] ), //i
    .b   (dSP_1038_b[7:0] ), //i
    .p   (dSP_1038_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1039 (
    .a   (dSP_1039_a[7:0] ), //i
    .d   (dSP_1039_d[7:0] ), //i
    .b   (dSP_1039_b[7:0] ), //i
    .p   (dSP_1039_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1040 (
    .a   (dSP_1040_a[7:0] ), //i
    .d   (dSP_1040_d[7:0] ), //i
    .b   (dSP_1040_b[7:0] ), //i
    .p   (dSP_1040_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1041 (
    .a   (dSP_1041_a[7:0] ), //i
    .d   (dSP_1041_d[7:0] ), //i
    .b   (dSP_1041_b[7:0] ), //i
    .p   (dSP_1041_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1042 (
    .a   (dSP_1042_a[7:0] ), //i
    .d   (dSP_1042_d[7:0] ), //i
    .b   (dSP_1042_b[7:0] ), //i
    .p   (dSP_1042_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1043 (
    .a   (dSP_1043_a[7:0] ), //i
    .d   (dSP_1043_d[7:0] ), //i
    .b   (dSP_1043_b[7:0] ), //i
    .p   (dSP_1043_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1044 (
    .a   (dSP_1044_a[7:0] ), //i
    .d   (dSP_1044_d[7:0] ), //i
    .b   (dSP_1044_b[7:0] ), //i
    .p   (dSP_1044_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1045 (
    .a   (dSP_1045_a[7:0] ), //i
    .d   (dSP_1045_d[7:0] ), //i
    .b   (dSP_1045_b[7:0] ), //i
    .p   (dSP_1045_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1046 (
    .a   (dSP_1046_a[7:0] ), //i
    .d   (dSP_1046_d[7:0] ), //i
    .b   (dSP_1046_b[7:0] ), //i
    .p   (dSP_1046_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1047 (
    .a   (dSP_1047_a[7:0] ), //i
    .d   (dSP_1047_d[7:0] ), //i
    .b   (dSP_1047_b[7:0] ), //i
    .p   (dSP_1047_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1048 (
    .a   (dSP_1048_a[7:0] ), //i
    .d   (dSP_1048_d[7:0] ), //i
    .b   (dSP_1048_b[7:0] ), //i
    .p   (dSP_1048_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1049 (
    .a   (dSP_1049_a[7:0] ), //i
    .d   (dSP_1049_d[7:0] ), //i
    .b   (dSP_1049_b[7:0] ), //i
    .p   (dSP_1049_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1050 (
    .a   (dSP_1050_a[7:0] ), //i
    .d   (dSP_1050_d[7:0] ), //i
    .b   (dSP_1050_b[7:0] ), //i
    .p   (dSP_1050_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1051 (
    .a   (dSP_1051_a[7:0] ), //i
    .d   (dSP_1051_d[7:0] ), //i
    .b   (dSP_1051_b[7:0] ), //i
    .p   (dSP_1051_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1052 (
    .a   (dSP_1052_a[7:0] ), //i
    .d   (dSP_1052_d[7:0] ), //i
    .b   (dSP_1052_b[7:0] ), //i
    .p   (dSP_1052_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1053 (
    .a   (dSP_1053_a[7:0] ), //i
    .d   (dSP_1053_d[7:0] ), //i
    .b   (dSP_1053_b[7:0] ), //i
    .p   (dSP_1053_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1054 (
    .a   (dSP_1054_a[7:0] ), //i
    .d   (dSP_1054_d[7:0] ), //i
    .b   (dSP_1054_b[7:0] ), //i
    .p   (dSP_1054_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1055 (
    .a   (dSP_1055_a[7:0] ), //i
    .d   (dSP_1055_d[7:0] ), //i
    .b   (dSP_1055_b[7:0] ), //i
    .p   (dSP_1055_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1056 (
    .a   (dSP_1056_a[7:0] ), //i
    .d   (dSP_1056_d[7:0] ), //i
    .b   (dSP_1056_b[7:0] ), //i
    .p   (dSP_1056_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1057 (
    .a   (dSP_1057_a[7:0] ), //i
    .d   (dSP_1057_d[7:0] ), //i
    .b   (dSP_1057_b[7:0] ), //i
    .p   (dSP_1057_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1058 (
    .a   (dSP_1058_a[7:0] ), //i
    .d   (dSP_1058_d[7:0] ), //i
    .b   (dSP_1058_b[7:0] ), //i
    .p   (dSP_1058_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1059 (
    .a   (dSP_1059_a[7:0] ), //i
    .d   (dSP_1059_d[7:0] ), //i
    .b   (dSP_1059_b[7:0] ), //i
    .p   (dSP_1059_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1060 (
    .a   (dSP_1060_a[7:0] ), //i
    .d   (dSP_1060_d[7:0] ), //i
    .b   (dSP_1060_b[7:0] ), //i
    .p   (dSP_1060_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1061 (
    .a   (dSP_1061_a[7:0] ), //i
    .d   (dSP_1061_d[7:0] ), //i
    .b   (dSP_1061_b[7:0] ), //i
    .p   (dSP_1061_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1062 (
    .a   (dSP_1062_a[7:0] ), //i
    .d   (dSP_1062_d[7:0] ), //i
    .b   (dSP_1062_b[7:0] ), //i
    .p   (dSP_1062_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1063 (
    .a   (dSP_1063_a[7:0] ), //i
    .d   (dSP_1063_d[7:0] ), //i
    .b   (dSP_1063_b[7:0] ), //i
    .p   (dSP_1063_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1064 (
    .a   (dSP_1064_a[7:0] ), //i
    .d   (dSP_1064_d[7:0] ), //i
    .b   (dSP_1064_b[7:0] ), //i
    .p   (dSP_1064_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1065 (
    .a   (dSP_1065_a[7:0] ), //i
    .d   (dSP_1065_d[7:0] ), //i
    .b   (dSP_1065_b[7:0] ), //i
    .p   (dSP_1065_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1066 (
    .a   (dSP_1066_a[7:0] ), //i
    .d   (dSP_1066_d[7:0] ), //i
    .b   (dSP_1066_b[7:0] ), //i
    .p   (dSP_1066_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1067 (
    .a   (dSP_1067_a[7:0] ), //i
    .d   (dSP_1067_d[7:0] ), //i
    .b   (dSP_1067_b[7:0] ), //i
    .p   (dSP_1067_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1068 (
    .a   (dSP_1068_a[7:0] ), //i
    .d   (dSP_1068_d[7:0] ), //i
    .b   (dSP_1068_b[7:0] ), //i
    .p   (dSP_1068_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1069 (
    .a   (dSP_1069_a[7:0] ), //i
    .d   (dSP_1069_d[7:0] ), //i
    .b   (dSP_1069_b[7:0] ), //i
    .p   (dSP_1069_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1070 (
    .a   (dSP_1070_a[7:0] ), //i
    .d   (dSP_1070_d[7:0] ), //i
    .b   (dSP_1070_b[7:0] ), //i
    .p   (dSP_1070_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1071 (
    .a   (dSP_1071_a[7:0] ), //i
    .d   (dSP_1071_d[7:0] ), //i
    .b   (dSP_1071_b[7:0] ), //i
    .p   (dSP_1071_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1072 (
    .a   (dSP_1072_a[7:0] ), //i
    .d   (dSP_1072_d[7:0] ), //i
    .b   (dSP_1072_b[7:0] ), //i
    .p   (dSP_1072_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1073 (
    .a   (dSP_1073_a[7:0] ), //i
    .d   (dSP_1073_d[7:0] ), //i
    .b   (dSP_1073_b[7:0] ), //i
    .p   (dSP_1073_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1074 (
    .a   (dSP_1074_a[7:0] ), //i
    .d   (dSP_1074_d[7:0] ), //i
    .b   (dSP_1074_b[7:0] ), //i
    .p   (dSP_1074_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1075 (
    .a   (dSP_1075_a[7:0] ), //i
    .d   (dSP_1075_d[7:0] ), //i
    .b   (dSP_1075_b[7:0] ), //i
    .p   (dSP_1075_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1076 (
    .a   (dSP_1076_a[7:0] ), //i
    .d   (dSP_1076_d[7:0] ), //i
    .b   (dSP_1076_b[7:0] ), //i
    .p   (dSP_1076_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1077 (
    .a   (dSP_1077_a[7:0] ), //i
    .d   (dSP_1077_d[7:0] ), //i
    .b   (dSP_1077_b[7:0] ), //i
    .p   (dSP_1077_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1078 (
    .a   (dSP_1078_a[7:0] ), //i
    .d   (dSP_1078_d[7:0] ), //i
    .b   (dSP_1078_b[7:0] ), //i
    .p   (dSP_1078_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1079 (
    .a   (dSP_1079_a[7:0] ), //i
    .d   (dSP_1079_d[7:0] ), //i
    .b   (dSP_1079_b[7:0] ), //i
    .p   (dSP_1079_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1080 (
    .a   (dSP_1080_a[7:0] ), //i
    .d   (dSP_1080_d[7:0] ), //i
    .b   (dSP_1080_b[7:0] ), //i
    .p   (dSP_1080_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1081 (
    .a   (dSP_1081_a[7:0] ), //i
    .d   (dSP_1081_d[7:0] ), //i
    .b   (dSP_1081_b[7:0] ), //i
    .p   (dSP_1081_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1082 (
    .a   (dSP_1082_a[7:0] ), //i
    .d   (dSP_1082_d[7:0] ), //i
    .b   (dSP_1082_b[7:0] ), //i
    .p   (dSP_1082_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1083 (
    .a   (dSP_1083_a[7:0] ), //i
    .d   (dSP_1083_d[7:0] ), //i
    .b   (dSP_1083_b[7:0] ), //i
    .p   (dSP_1083_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1084 (
    .a   (dSP_1084_a[7:0] ), //i
    .d   (dSP_1084_d[7:0] ), //i
    .b   (dSP_1084_b[7:0] ), //i
    .p   (dSP_1084_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1085 (
    .a   (dSP_1085_a[7:0] ), //i
    .d   (dSP_1085_d[7:0] ), //i
    .b   (dSP_1085_b[7:0] ), //i
    .p   (dSP_1085_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1086 (
    .a   (dSP_1086_a[7:0] ), //i
    .d   (dSP_1086_d[7:0] ), //i
    .b   (dSP_1086_b[7:0] ), //i
    .p   (dSP_1086_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1087 (
    .a   (dSP_1087_a[7:0] ), //i
    .d   (dSP_1087_d[7:0] ), //i
    .b   (dSP_1087_b[7:0] ), //i
    .p   (dSP_1087_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1088 (
    .a   (dSP_1088_a[7:0] ), //i
    .d   (dSP_1088_d[7:0] ), //i
    .b   (dSP_1088_b[7:0] ), //i
    .p   (dSP_1088_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1089 (
    .a   (dSP_1089_a[7:0] ), //i
    .d   (dSP_1089_d[7:0] ), //i
    .b   (dSP_1089_b[7:0] ), //i
    .p   (dSP_1089_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1090 (
    .a   (dSP_1090_a[7:0] ), //i
    .d   (dSP_1090_d[7:0] ), //i
    .b   (dSP_1090_b[7:0] ), //i
    .p   (dSP_1090_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1091 (
    .a   (dSP_1091_a[7:0] ), //i
    .d   (dSP_1091_d[7:0] ), //i
    .b   (dSP_1091_b[7:0] ), //i
    .p   (dSP_1091_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1092 (
    .a   (dSP_1092_a[7:0] ), //i
    .d   (dSP_1092_d[7:0] ), //i
    .b   (dSP_1092_b[7:0] ), //i
    .p   (dSP_1092_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1093 (
    .a   (dSP_1093_a[7:0] ), //i
    .d   (dSP_1093_d[7:0] ), //i
    .b   (dSP_1093_b[7:0] ), //i
    .p   (dSP_1093_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1094 (
    .a   (dSP_1094_a[7:0] ), //i
    .d   (dSP_1094_d[7:0] ), //i
    .b   (dSP_1094_b[7:0] ), //i
    .p   (dSP_1094_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1095 (
    .a   (dSP_1095_a[7:0] ), //i
    .d   (dSP_1095_d[7:0] ), //i
    .b   (dSP_1095_b[7:0] ), //i
    .p   (dSP_1095_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1096 (
    .a   (dSP_1096_a[7:0] ), //i
    .d   (dSP_1096_d[7:0] ), //i
    .b   (dSP_1096_b[7:0] ), //i
    .p   (dSP_1096_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1097 (
    .a   (dSP_1097_a[7:0] ), //i
    .d   (dSP_1097_d[7:0] ), //i
    .b   (dSP_1097_b[7:0] ), //i
    .p   (dSP_1097_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1098 (
    .a   (dSP_1098_a[7:0] ), //i
    .d   (dSP_1098_d[7:0] ), //i
    .b   (dSP_1098_b[7:0] ), //i
    .p   (dSP_1098_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1099 (
    .a   (dSP_1099_a[7:0] ), //i
    .d   (dSP_1099_d[7:0] ), //i
    .b   (dSP_1099_b[7:0] ), //i
    .p   (dSP_1099_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1100 (
    .a   (dSP_1100_a[7:0] ), //i
    .d   (dSP_1100_d[7:0] ), //i
    .b   (dSP_1100_b[7:0] ), //i
    .p   (dSP_1100_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1101 (
    .a   (dSP_1101_a[7:0] ), //i
    .d   (dSP_1101_d[7:0] ), //i
    .b   (dSP_1101_b[7:0] ), //i
    .p   (dSP_1101_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1102 (
    .a   (dSP_1102_a[7:0] ), //i
    .d   (dSP_1102_d[7:0] ), //i
    .b   (dSP_1102_b[7:0] ), //i
    .p   (dSP_1102_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1103 (
    .a   (dSP_1103_a[7:0] ), //i
    .d   (dSP_1103_d[7:0] ), //i
    .b   (dSP_1103_b[7:0] ), //i
    .p   (dSP_1103_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1104 (
    .a   (dSP_1104_a[7:0] ), //i
    .d   (dSP_1104_d[7:0] ), //i
    .b   (dSP_1104_b[7:0] ), //i
    .p   (dSP_1104_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1105 (
    .a   (dSP_1105_a[7:0] ), //i
    .d   (dSP_1105_d[7:0] ), //i
    .b   (dSP_1105_b[7:0] ), //i
    .p   (dSP_1105_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1106 (
    .a   (dSP_1106_a[7:0] ), //i
    .d   (dSP_1106_d[7:0] ), //i
    .b   (dSP_1106_b[7:0] ), //i
    .p   (dSP_1106_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1107 (
    .a   (dSP_1107_a[7:0] ), //i
    .d   (dSP_1107_d[7:0] ), //i
    .b   (dSP_1107_b[7:0] ), //i
    .p   (dSP_1107_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1108 (
    .a   (dSP_1108_a[7:0] ), //i
    .d   (dSP_1108_d[7:0] ), //i
    .b   (dSP_1108_b[7:0] ), //i
    .p   (dSP_1108_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1109 (
    .a   (dSP_1109_a[7:0] ), //i
    .d   (dSP_1109_d[7:0] ), //i
    .b   (dSP_1109_b[7:0] ), //i
    .p   (dSP_1109_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1110 (
    .a   (dSP_1110_a[7:0] ), //i
    .d   (dSP_1110_d[7:0] ), //i
    .b   (dSP_1110_b[7:0] ), //i
    .p   (dSP_1110_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1111 (
    .a   (dSP_1111_a[7:0] ), //i
    .d   (dSP_1111_d[7:0] ), //i
    .b   (dSP_1111_b[7:0] ), //i
    .p   (dSP_1111_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1112 (
    .a   (dSP_1112_a[7:0] ), //i
    .d   (dSP_1112_d[7:0] ), //i
    .b   (dSP_1112_b[7:0] ), //i
    .p   (dSP_1112_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1113 (
    .a   (dSP_1113_a[7:0] ), //i
    .d   (dSP_1113_d[7:0] ), //i
    .b   (dSP_1113_b[7:0] ), //i
    .p   (dSP_1113_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1114 (
    .a   (dSP_1114_a[7:0] ), //i
    .d   (dSP_1114_d[7:0] ), //i
    .b   (dSP_1114_b[7:0] ), //i
    .p   (dSP_1114_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1115 (
    .a   (dSP_1115_a[7:0] ), //i
    .d   (dSP_1115_d[7:0] ), //i
    .b   (dSP_1115_b[7:0] ), //i
    .p   (dSP_1115_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1116 (
    .a   (dSP_1116_a[7:0] ), //i
    .d   (dSP_1116_d[7:0] ), //i
    .b   (dSP_1116_b[7:0] ), //i
    .p   (dSP_1116_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1117 (
    .a   (dSP_1117_a[7:0] ), //i
    .d   (dSP_1117_d[7:0] ), //i
    .b   (dSP_1117_b[7:0] ), //i
    .p   (dSP_1117_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1118 (
    .a   (dSP_1118_a[7:0] ), //i
    .d   (dSP_1118_d[7:0] ), //i
    .b   (dSP_1118_b[7:0] ), //i
    .p   (dSP_1118_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1119 (
    .a   (dSP_1119_a[7:0] ), //i
    .d   (dSP_1119_d[7:0] ), //i
    .b   (dSP_1119_b[7:0] ), //i
    .p   (dSP_1119_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1120 (
    .a   (dSP_1120_a[7:0] ), //i
    .d   (dSP_1120_d[7:0] ), //i
    .b   (dSP_1120_b[7:0] ), //i
    .p   (dSP_1120_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1121 (
    .a   (dSP_1121_a[7:0] ), //i
    .d   (dSP_1121_d[7:0] ), //i
    .b   (dSP_1121_b[7:0] ), //i
    .p   (dSP_1121_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1122 (
    .a   (dSP_1122_a[7:0] ), //i
    .d   (dSP_1122_d[7:0] ), //i
    .b   (dSP_1122_b[7:0] ), //i
    .p   (dSP_1122_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1123 (
    .a   (dSP_1123_a[7:0] ), //i
    .d   (dSP_1123_d[7:0] ), //i
    .b   (dSP_1123_b[7:0] ), //i
    .p   (dSP_1123_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1124 (
    .a   (dSP_1124_a[7:0] ), //i
    .d   (dSP_1124_d[7:0] ), //i
    .b   (dSP_1124_b[7:0] ), //i
    .p   (dSP_1124_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1125 (
    .a   (dSP_1125_a[7:0] ), //i
    .d   (dSP_1125_d[7:0] ), //i
    .b   (dSP_1125_b[7:0] ), //i
    .p   (dSP_1125_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1126 (
    .a   (dSP_1126_a[7:0] ), //i
    .d   (dSP_1126_d[7:0] ), //i
    .b   (dSP_1126_b[7:0] ), //i
    .p   (dSP_1126_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1127 (
    .a   (dSP_1127_a[7:0] ), //i
    .d   (dSP_1127_d[7:0] ), //i
    .b   (dSP_1127_b[7:0] ), //i
    .p   (dSP_1127_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1128 (
    .a   (dSP_1128_a[7:0] ), //i
    .d   (dSP_1128_d[7:0] ), //i
    .b   (dSP_1128_b[7:0] ), //i
    .p   (dSP_1128_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1129 (
    .a   (dSP_1129_a[7:0] ), //i
    .d   (dSP_1129_d[7:0] ), //i
    .b   (dSP_1129_b[7:0] ), //i
    .p   (dSP_1129_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1130 (
    .a   (dSP_1130_a[7:0] ), //i
    .d   (dSP_1130_d[7:0] ), //i
    .b   (dSP_1130_b[7:0] ), //i
    .p   (dSP_1130_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1131 (
    .a   (dSP_1131_a[7:0] ), //i
    .d   (dSP_1131_d[7:0] ), //i
    .b   (dSP_1131_b[7:0] ), //i
    .p   (dSP_1131_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1132 (
    .a   (dSP_1132_a[7:0] ), //i
    .d   (dSP_1132_d[7:0] ), //i
    .b   (dSP_1132_b[7:0] ), //i
    .p   (dSP_1132_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1133 (
    .a   (dSP_1133_a[7:0] ), //i
    .d   (dSP_1133_d[7:0] ), //i
    .b   (dSP_1133_b[7:0] ), //i
    .p   (dSP_1133_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1134 (
    .a   (dSP_1134_a[7:0] ), //i
    .d   (dSP_1134_d[7:0] ), //i
    .b   (dSP_1134_b[7:0] ), //i
    .p   (dSP_1134_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1135 (
    .a   (dSP_1135_a[7:0] ), //i
    .d   (dSP_1135_d[7:0] ), //i
    .b   (dSP_1135_b[7:0] ), //i
    .p   (dSP_1135_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1136 (
    .a   (dSP_1136_a[7:0] ), //i
    .d   (dSP_1136_d[7:0] ), //i
    .b   (dSP_1136_b[7:0] ), //i
    .p   (dSP_1136_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1137 (
    .a   (dSP_1137_a[7:0] ), //i
    .d   (dSP_1137_d[7:0] ), //i
    .b   (dSP_1137_b[7:0] ), //i
    .p   (dSP_1137_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1138 (
    .a   (dSP_1138_a[7:0] ), //i
    .d   (dSP_1138_d[7:0] ), //i
    .b   (dSP_1138_b[7:0] ), //i
    .p   (dSP_1138_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1139 (
    .a   (dSP_1139_a[7:0] ), //i
    .d   (dSP_1139_d[7:0] ), //i
    .b   (dSP_1139_b[7:0] ), //i
    .p   (dSP_1139_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1140 (
    .a   (dSP_1140_a[7:0] ), //i
    .d   (dSP_1140_d[7:0] ), //i
    .b   (dSP_1140_b[7:0] ), //i
    .p   (dSP_1140_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1141 (
    .a   (dSP_1141_a[7:0] ), //i
    .d   (dSP_1141_d[7:0] ), //i
    .b   (dSP_1141_b[7:0] ), //i
    .p   (dSP_1141_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1142 (
    .a   (dSP_1142_a[7:0] ), //i
    .d   (dSP_1142_d[7:0] ), //i
    .b   (dSP_1142_b[7:0] ), //i
    .p   (dSP_1142_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1143 (
    .a   (dSP_1143_a[7:0] ), //i
    .d   (dSP_1143_d[7:0] ), //i
    .b   (dSP_1143_b[7:0] ), //i
    .p   (dSP_1143_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1144 (
    .a   (dSP_1144_a[7:0] ), //i
    .d   (dSP_1144_d[7:0] ), //i
    .b   (dSP_1144_b[7:0] ), //i
    .p   (dSP_1144_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1145 (
    .a   (dSP_1145_a[7:0] ), //i
    .d   (dSP_1145_d[7:0] ), //i
    .b   (dSP_1145_b[7:0] ), //i
    .p   (dSP_1145_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1146 (
    .a   (dSP_1146_a[7:0] ), //i
    .d   (dSP_1146_d[7:0] ), //i
    .b   (dSP_1146_b[7:0] ), //i
    .p   (dSP_1146_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1147 (
    .a   (dSP_1147_a[7:0] ), //i
    .d   (dSP_1147_d[7:0] ), //i
    .b   (dSP_1147_b[7:0] ), //i
    .p   (dSP_1147_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1148 (
    .a   (dSP_1148_a[7:0] ), //i
    .d   (dSP_1148_d[7:0] ), //i
    .b   (dSP_1148_b[7:0] ), //i
    .p   (dSP_1148_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1149 (
    .a   (dSP_1149_a[7:0] ), //i
    .d   (dSP_1149_d[7:0] ), //i
    .b   (dSP_1149_b[7:0] ), //i
    .p   (dSP_1149_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1150 (
    .a   (dSP_1150_a[7:0] ), //i
    .d   (dSP_1150_d[7:0] ), //i
    .b   (dSP_1150_b[7:0] ), //i
    .p   (dSP_1150_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1151 (
    .a   (dSP_1151_a[7:0] ), //i
    .d   (dSP_1151_d[7:0] ), //i
    .b   (dSP_1151_b[7:0] ), //i
    .p   (dSP_1151_p[31:0]), //o
    .CLK (clk             )  //i
  );
  DSP dSP_1152 (
    .a   (dSP_1152_a[7:0] ), //i
    .d   (dSP_1152_d[7:0] ), //i
    .b   (dSP_1152_b[7:0] ), //i
    .p   (dSP_1152_p[31:0]), //o
    .CLK (clk             )  //i
  );
  xAddTimes addKernel (
    .A_0       (addKernel_A_0[31:0]), //i
    .A_1       (addKernel_A_1[31:0]), //i
    .A_2       (addKernel_A_2[31:0]), //i
    .A_3       (addKernel_A_3[31:0]), //i
    .A_4       (addKernel_A_4[31:0]), //i
    .A_5       (addKernel_A_5[31:0]), //i
    .A_6       (addKernel_A_6[31:0]), //i
    .A_7       (addKernel_A_7[31:0]), //i
    .A_8       (addKernel_A_8[31:0]), //i
    .S         (addKernel_S[39:0]  ), //o
    .clk       (clk                ), //i
    .reset     (reset              ), //i
    .softReset (softReset          )  //i
  );
  xAddTimes addKernel_1 (
    .A_0       (addKernel_1_A_0[31:0]), //i
    .A_1       (addKernel_1_A_1[31:0]), //i
    .A_2       (addKernel_1_A_2[31:0]), //i
    .A_3       (addKernel_1_A_3[31:0]), //i
    .A_4       (addKernel_1_A_4[31:0]), //i
    .A_5       (addKernel_1_A_5[31:0]), //i
    .A_6       (addKernel_1_A_6[31:0]), //i
    .A_7       (addKernel_1_A_7[31:0]), //i
    .A_8       (addKernel_1_A_8[31:0]), //i
    .S         (addKernel_1_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_2 (
    .A_0       (addKernel_2_A_0[31:0]), //i
    .A_1       (addKernel_2_A_1[31:0]), //i
    .A_2       (addKernel_2_A_2[31:0]), //i
    .A_3       (addKernel_2_A_3[31:0]), //i
    .A_4       (addKernel_2_A_4[31:0]), //i
    .A_5       (addKernel_2_A_5[31:0]), //i
    .A_6       (addKernel_2_A_6[31:0]), //i
    .A_7       (addKernel_2_A_7[31:0]), //i
    .A_8       (addKernel_2_A_8[31:0]), //i
    .S         (addKernel_2_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_3 (
    .A_0       (addKernel_3_A_0[31:0]), //i
    .A_1       (addKernel_3_A_1[31:0]), //i
    .A_2       (addKernel_3_A_2[31:0]), //i
    .A_3       (addKernel_3_A_3[31:0]), //i
    .A_4       (addKernel_3_A_4[31:0]), //i
    .A_5       (addKernel_3_A_5[31:0]), //i
    .A_6       (addKernel_3_A_6[31:0]), //i
    .A_7       (addKernel_3_A_7[31:0]), //i
    .A_8       (addKernel_3_A_8[31:0]), //i
    .S         (addKernel_3_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_4 (
    .A_0       (addKernel_4_A_0[31:0]), //i
    .A_1       (addKernel_4_A_1[31:0]), //i
    .A_2       (addKernel_4_A_2[31:0]), //i
    .A_3       (addKernel_4_A_3[31:0]), //i
    .A_4       (addKernel_4_A_4[31:0]), //i
    .A_5       (addKernel_4_A_5[31:0]), //i
    .A_6       (addKernel_4_A_6[31:0]), //i
    .A_7       (addKernel_4_A_7[31:0]), //i
    .A_8       (addKernel_4_A_8[31:0]), //i
    .S         (addKernel_4_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_5 (
    .A_0       (addKernel_5_A_0[31:0]), //i
    .A_1       (addKernel_5_A_1[31:0]), //i
    .A_2       (addKernel_5_A_2[31:0]), //i
    .A_3       (addKernel_5_A_3[31:0]), //i
    .A_4       (addKernel_5_A_4[31:0]), //i
    .A_5       (addKernel_5_A_5[31:0]), //i
    .A_6       (addKernel_5_A_6[31:0]), //i
    .A_7       (addKernel_5_A_7[31:0]), //i
    .A_8       (addKernel_5_A_8[31:0]), //i
    .S         (addKernel_5_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_6 (
    .A_0       (addKernel_6_A_0[31:0]), //i
    .A_1       (addKernel_6_A_1[31:0]), //i
    .A_2       (addKernel_6_A_2[31:0]), //i
    .A_3       (addKernel_6_A_3[31:0]), //i
    .A_4       (addKernel_6_A_4[31:0]), //i
    .A_5       (addKernel_6_A_5[31:0]), //i
    .A_6       (addKernel_6_A_6[31:0]), //i
    .A_7       (addKernel_6_A_7[31:0]), //i
    .A_8       (addKernel_6_A_8[31:0]), //i
    .S         (addKernel_6_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_7 (
    .A_0       (addKernel_7_A_0[31:0]), //i
    .A_1       (addKernel_7_A_1[31:0]), //i
    .A_2       (addKernel_7_A_2[31:0]), //i
    .A_3       (addKernel_7_A_3[31:0]), //i
    .A_4       (addKernel_7_A_4[31:0]), //i
    .A_5       (addKernel_7_A_5[31:0]), //i
    .A_6       (addKernel_7_A_6[31:0]), //i
    .A_7       (addKernel_7_A_7[31:0]), //i
    .A_8       (addKernel_7_A_8[31:0]), //i
    .S         (addKernel_7_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_8 (
    .A_0       (addKernel_8_A_0[31:0]), //i
    .A_1       (addKernel_8_A_1[31:0]), //i
    .A_2       (addKernel_8_A_2[31:0]), //i
    .A_3       (addKernel_8_A_3[31:0]), //i
    .A_4       (addKernel_8_A_4[31:0]), //i
    .A_5       (addKernel_8_A_5[31:0]), //i
    .A_6       (addKernel_8_A_6[31:0]), //i
    .A_7       (addKernel_8_A_7[31:0]), //i
    .A_8       (addKernel_8_A_8[31:0]), //i
    .S         (addKernel_8_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_9 (
    .A_0       (addKernel_9_A_0[31:0]), //i
    .A_1       (addKernel_9_A_1[31:0]), //i
    .A_2       (addKernel_9_A_2[31:0]), //i
    .A_3       (addKernel_9_A_3[31:0]), //i
    .A_4       (addKernel_9_A_4[31:0]), //i
    .A_5       (addKernel_9_A_5[31:0]), //i
    .A_6       (addKernel_9_A_6[31:0]), //i
    .A_7       (addKernel_9_A_7[31:0]), //i
    .A_8       (addKernel_9_A_8[31:0]), //i
    .S         (addKernel_9_S[39:0]  ), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes addKernel_10 (
    .A_0       (addKernel_10_A_0[31:0]), //i
    .A_1       (addKernel_10_A_1[31:0]), //i
    .A_2       (addKernel_10_A_2[31:0]), //i
    .A_3       (addKernel_10_A_3[31:0]), //i
    .A_4       (addKernel_10_A_4[31:0]), //i
    .A_5       (addKernel_10_A_5[31:0]), //i
    .A_6       (addKernel_10_A_6[31:0]), //i
    .A_7       (addKernel_10_A_7[31:0]), //i
    .A_8       (addKernel_10_A_8[31:0]), //i
    .S         (addKernel_10_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_11 (
    .A_0       (addKernel_11_A_0[31:0]), //i
    .A_1       (addKernel_11_A_1[31:0]), //i
    .A_2       (addKernel_11_A_2[31:0]), //i
    .A_3       (addKernel_11_A_3[31:0]), //i
    .A_4       (addKernel_11_A_4[31:0]), //i
    .A_5       (addKernel_11_A_5[31:0]), //i
    .A_6       (addKernel_11_A_6[31:0]), //i
    .A_7       (addKernel_11_A_7[31:0]), //i
    .A_8       (addKernel_11_A_8[31:0]), //i
    .S         (addKernel_11_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_12 (
    .A_0       (addKernel_12_A_0[31:0]), //i
    .A_1       (addKernel_12_A_1[31:0]), //i
    .A_2       (addKernel_12_A_2[31:0]), //i
    .A_3       (addKernel_12_A_3[31:0]), //i
    .A_4       (addKernel_12_A_4[31:0]), //i
    .A_5       (addKernel_12_A_5[31:0]), //i
    .A_6       (addKernel_12_A_6[31:0]), //i
    .A_7       (addKernel_12_A_7[31:0]), //i
    .A_8       (addKernel_12_A_8[31:0]), //i
    .S         (addKernel_12_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_13 (
    .A_0       (addKernel_13_A_0[31:0]), //i
    .A_1       (addKernel_13_A_1[31:0]), //i
    .A_2       (addKernel_13_A_2[31:0]), //i
    .A_3       (addKernel_13_A_3[31:0]), //i
    .A_4       (addKernel_13_A_4[31:0]), //i
    .A_5       (addKernel_13_A_5[31:0]), //i
    .A_6       (addKernel_13_A_6[31:0]), //i
    .A_7       (addKernel_13_A_7[31:0]), //i
    .A_8       (addKernel_13_A_8[31:0]), //i
    .S         (addKernel_13_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_14 (
    .A_0       (addKernel_14_A_0[31:0]), //i
    .A_1       (addKernel_14_A_1[31:0]), //i
    .A_2       (addKernel_14_A_2[31:0]), //i
    .A_3       (addKernel_14_A_3[31:0]), //i
    .A_4       (addKernel_14_A_4[31:0]), //i
    .A_5       (addKernel_14_A_5[31:0]), //i
    .A_6       (addKernel_14_A_6[31:0]), //i
    .A_7       (addKernel_14_A_7[31:0]), //i
    .A_8       (addKernel_14_A_8[31:0]), //i
    .S         (addKernel_14_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_15 (
    .A_0       (addKernel_15_A_0[31:0]), //i
    .A_1       (addKernel_15_A_1[31:0]), //i
    .A_2       (addKernel_15_A_2[31:0]), //i
    .A_3       (addKernel_15_A_3[31:0]), //i
    .A_4       (addKernel_15_A_4[31:0]), //i
    .A_5       (addKernel_15_A_5[31:0]), //i
    .A_6       (addKernel_15_A_6[31:0]), //i
    .A_7       (addKernel_15_A_7[31:0]), //i
    .A_8       (addKernel_15_A_8[31:0]), //i
    .S         (addKernel_15_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_16 (
    .A_0       (addKernel_16_A_0[31:0]), //i
    .A_1       (addKernel_16_A_1[31:0]), //i
    .A_2       (addKernel_16_A_2[31:0]), //i
    .A_3       (addKernel_16_A_3[31:0]), //i
    .A_4       (addKernel_16_A_4[31:0]), //i
    .A_5       (addKernel_16_A_5[31:0]), //i
    .A_6       (addKernel_16_A_6[31:0]), //i
    .A_7       (addKernel_16_A_7[31:0]), //i
    .A_8       (addKernel_16_A_8[31:0]), //i
    .S         (addKernel_16_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_17 (
    .A_0       (addKernel_17_A_0[31:0]), //i
    .A_1       (addKernel_17_A_1[31:0]), //i
    .A_2       (addKernel_17_A_2[31:0]), //i
    .A_3       (addKernel_17_A_3[31:0]), //i
    .A_4       (addKernel_17_A_4[31:0]), //i
    .A_5       (addKernel_17_A_5[31:0]), //i
    .A_6       (addKernel_17_A_6[31:0]), //i
    .A_7       (addKernel_17_A_7[31:0]), //i
    .A_8       (addKernel_17_A_8[31:0]), //i
    .S         (addKernel_17_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_18 (
    .A_0       (addKernel_18_A_0[31:0]), //i
    .A_1       (addKernel_18_A_1[31:0]), //i
    .A_2       (addKernel_18_A_2[31:0]), //i
    .A_3       (addKernel_18_A_3[31:0]), //i
    .A_4       (addKernel_18_A_4[31:0]), //i
    .A_5       (addKernel_18_A_5[31:0]), //i
    .A_6       (addKernel_18_A_6[31:0]), //i
    .A_7       (addKernel_18_A_7[31:0]), //i
    .A_8       (addKernel_18_A_8[31:0]), //i
    .S         (addKernel_18_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_19 (
    .A_0       (addKernel_19_A_0[31:0]), //i
    .A_1       (addKernel_19_A_1[31:0]), //i
    .A_2       (addKernel_19_A_2[31:0]), //i
    .A_3       (addKernel_19_A_3[31:0]), //i
    .A_4       (addKernel_19_A_4[31:0]), //i
    .A_5       (addKernel_19_A_5[31:0]), //i
    .A_6       (addKernel_19_A_6[31:0]), //i
    .A_7       (addKernel_19_A_7[31:0]), //i
    .A_8       (addKernel_19_A_8[31:0]), //i
    .S         (addKernel_19_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_20 (
    .A_0       (addKernel_20_A_0[31:0]), //i
    .A_1       (addKernel_20_A_1[31:0]), //i
    .A_2       (addKernel_20_A_2[31:0]), //i
    .A_3       (addKernel_20_A_3[31:0]), //i
    .A_4       (addKernel_20_A_4[31:0]), //i
    .A_5       (addKernel_20_A_5[31:0]), //i
    .A_6       (addKernel_20_A_6[31:0]), //i
    .A_7       (addKernel_20_A_7[31:0]), //i
    .A_8       (addKernel_20_A_8[31:0]), //i
    .S         (addKernel_20_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_21 (
    .A_0       (addKernel_21_A_0[31:0]), //i
    .A_1       (addKernel_21_A_1[31:0]), //i
    .A_2       (addKernel_21_A_2[31:0]), //i
    .A_3       (addKernel_21_A_3[31:0]), //i
    .A_4       (addKernel_21_A_4[31:0]), //i
    .A_5       (addKernel_21_A_5[31:0]), //i
    .A_6       (addKernel_21_A_6[31:0]), //i
    .A_7       (addKernel_21_A_7[31:0]), //i
    .A_8       (addKernel_21_A_8[31:0]), //i
    .S         (addKernel_21_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_22 (
    .A_0       (addKernel_22_A_0[31:0]), //i
    .A_1       (addKernel_22_A_1[31:0]), //i
    .A_2       (addKernel_22_A_2[31:0]), //i
    .A_3       (addKernel_22_A_3[31:0]), //i
    .A_4       (addKernel_22_A_4[31:0]), //i
    .A_5       (addKernel_22_A_5[31:0]), //i
    .A_6       (addKernel_22_A_6[31:0]), //i
    .A_7       (addKernel_22_A_7[31:0]), //i
    .A_8       (addKernel_22_A_8[31:0]), //i
    .S         (addKernel_22_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_23 (
    .A_0       (addKernel_23_A_0[31:0]), //i
    .A_1       (addKernel_23_A_1[31:0]), //i
    .A_2       (addKernel_23_A_2[31:0]), //i
    .A_3       (addKernel_23_A_3[31:0]), //i
    .A_4       (addKernel_23_A_4[31:0]), //i
    .A_5       (addKernel_23_A_5[31:0]), //i
    .A_6       (addKernel_23_A_6[31:0]), //i
    .A_7       (addKernel_23_A_7[31:0]), //i
    .A_8       (addKernel_23_A_8[31:0]), //i
    .S         (addKernel_23_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_24 (
    .A_0       (addKernel_24_A_0[31:0]), //i
    .A_1       (addKernel_24_A_1[31:0]), //i
    .A_2       (addKernel_24_A_2[31:0]), //i
    .A_3       (addKernel_24_A_3[31:0]), //i
    .A_4       (addKernel_24_A_4[31:0]), //i
    .A_5       (addKernel_24_A_5[31:0]), //i
    .A_6       (addKernel_24_A_6[31:0]), //i
    .A_7       (addKernel_24_A_7[31:0]), //i
    .A_8       (addKernel_24_A_8[31:0]), //i
    .S         (addKernel_24_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_25 (
    .A_0       (addKernel_25_A_0[31:0]), //i
    .A_1       (addKernel_25_A_1[31:0]), //i
    .A_2       (addKernel_25_A_2[31:0]), //i
    .A_3       (addKernel_25_A_3[31:0]), //i
    .A_4       (addKernel_25_A_4[31:0]), //i
    .A_5       (addKernel_25_A_5[31:0]), //i
    .A_6       (addKernel_25_A_6[31:0]), //i
    .A_7       (addKernel_25_A_7[31:0]), //i
    .A_8       (addKernel_25_A_8[31:0]), //i
    .S         (addKernel_25_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_26 (
    .A_0       (addKernel_26_A_0[31:0]), //i
    .A_1       (addKernel_26_A_1[31:0]), //i
    .A_2       (addKernel_26_A_2[31:0]), //i
    .A_3       (addKernel_26_A_3[31:0]), //i
    .A_4       (addKernel_26_A_4[31:0]), //i
    .A_5       (addKernel_26_A_5[31:0]), //i
    .A_6       (addKernel_26_A_6[31:0]), //i
    .A_7       (addKernel_26_A_7[31:0]), //i
    .A_8       (addKernel_26_A_8[31:0]), //i
    .S         (addKernel_26_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_27 (
    .A_0       (addKernel_27_A_0[31:0]), //i
    .A_1       (addKernel_27_A_1[31:0]), //i
    .A_2       (addKernel_27_A_2[31:0]), //i
    .A_3       (addKernel_27_A_3[31:0]), //i
    .A_4       (addKernel_27_A_4[31:0]), //i
    .A_5       (addKernel_27_A_5[31:0]), //i
    .A_6       (addKernel_27_A_6[31:0]), //i
    .A_7       (addKernel_27_A_7[31:0]), //i
    .A_8       (addKernel_27_A_8[31:0]), //i
    .S         (addKernel_27_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_28 (
    .A_0       (addKernel_28_A_0[31:0]), //i
    .A_1       (addKernel_28_A_1[31:0]), //i
    .A_2       (addKernel_28_A_2[31:0]), //i
    .A_3       (addKernel_28_A_3[31:0]), //i
    .A_4       (addKernel_28_A_4[31:0]), //i
    .A_5       (addKernel_28_A_5[31:0]), //i
    .A_6       (addKernel_28_A_6[31:0]), //i
    .A_7       (addKernel_28_A_7[31:0]), //i
    .A_8       (addKernel_28_A_8[31:0]), //i
    .S         (addKernel_28_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_29 (
    .A_0       (addKernel_29_A_0[31:0]), //i
    .A_1       (addKernel_29_A_1[31:0]), //i
    .A_2       (addKernel_29_A_2[31:0]), //i
    .A_3       (addKernel_29_A_3[31:0]), //i
    .A_4       (addKernel_29_A_4[31:0]), //i
    .A_5       (addKernel_29_A_5[31:0]), //i
    .A_6       (addKernel_29_A_6[31:0]), //i
    .A_7       (addKernel_29_A_7[31:0]), //i
    .A_8       (addKernel_29_A_8[31:0]), //i
    .S         (addKernel_29_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_30 (
    .A_0       (addKernel_30_A_0[31:0]), //i
    .A_1       (addKernel_30_A_1[31:0]), //i
    .A_2       (addKernel_30_A_2[31:0]), //i
    .A_3       (addKernel_30_A_3[31:0]), //i
    .A_4       (addKernel_30_A_4[31:0]), //i
    .A_5       (addKernel_30_A_5[31:0]), //i
    .A_6       (addKernel_30_A_6[31:0]), //i
    .A_7       (addKernel_30_A_7[31:0]), //i
    .A_8       (addKernel_30_A_8[31:0]), //i
    .S         (addKernel_30_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_31 (
    .A_0       (addKernel_31_A_0[31:0]), //i
    .A_1       (addKernel_31_A_1[31:0]), //i
    .A_2       (addKernel_31_A_2[31:0]), //i
    .A_3       (addKernel_31_A_3[31:0]), //i
    .A_4       (addKernel_31_A_4[31:0]), //i
    .A_5       (addKernel_31_A_5[31:0]), //i
    .A_6       (addKernel_31_A_6[31:0]), //i
    .A_7       (addKernel_31_A_7[31:0]), //i
    .A_8       (addKernel_31_A_8[31:0]), //i
    .S         (addKernel_31_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_32 (
    .A_0       (addKernel_32_A_0[31:0]), //i
    .A_1       (addKernel_32_A_1[31:0]), //i
    .A_2       (addKernel_32_A_2[31:0]), //i
    .A_3       (addKernel_32_A_3[31:0]), //i
    .A_4       (addKernel_32_A_4[31:0]), //i
    .A_5       (addKernel_32_A_5[31:0]), //i
    .A_6       (addKernel_32_A_6[31:0]), //i
    .A_7       (addKernel_32_A_7[31:0]), //i
    .A_8       (addKernel_32_A_8[31:0]), //i
    .S         (addKernel_32_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_33 (
    .A_0       (addKernel_33_A_0[31:0]), //i
    .A_1       (addKernel_33_A_1[31:0]), //i
    .A_2       (addKernel_33_A_2[31:0]), //i
    .A_3       (addKernel_33_A_3[31:0]), //i
    .A_4       (addKernel_33_A_4[31:0]), //i
    .A_5       (addKernel_33_A_5[31:0]), //i
    .A_6       (addKernel_33_A_6[31:0]), //i
    .A_7       (addKernel_33_A_7[31:0]), //i
    .A_8       (addKernel_33_A_8[31:0]), //i
    .S         (addKernel_33_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_34 (
    .A_0       (addKernel_34_A_0[31:0]), //i
    .A_1       (addKernel_34_A_1[31:0]), //i
    .A_2       (addKernel_34_A_2[31:0]), //i
    .A_3       (addKernel_34_A_3[31:0]), //i
    .A_4       (addKernel_34_A_4[31:0]), //i
    .A_5       (addKernel_34_A_5[31:0]), //i
    .A_6       (addKernel_34_A_6[31:0]), //i
    .A_7       (addKernel_34_A_7[31:0]), //i
    .A_8       (addKernel_34_A_8[31:0]), //i
    .S         (addKernel_34_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_35 (
    .A_0       (addKernel_35_A_0[31:0]), //i
    .A_1       (addKernel_35_A_1[31:0]), //i
    .A_2       (addKernel_35_A_2[31:0]), //i
    .A_3       (addKernel_35_A_3[31:0]), //i
    .A_4       (addKernel_35_A_4[31:0]), //i
    .A_5       (addKernel_35_A_5[31:0]), //i
    .A_6       (addKernel_35_A_6[31:0]), //i
    .A_7       (addKernel_35_A_7[31:0]), //i
    .A_8       (addKernel_35_A_8[31:0]), //i
    .S         (addKernel_35_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_36 (
    .A_0       (addKernel_36_A_0[31:0]), //i
    .A_1       (addKernel_36_A_1[31:0]), //i
    .A_2       (addKernel_36_A_2[31:0]), //i
    .A_3       (addKernel_36_A_3[31:0]), //i
    .A_4       (addKernel_36_A_4[31:0]), //i
    .A_5       (addKernel_36_A_5[31:0]), //i
    .A_6       (addKernel_36_A_6[31:0]), //i
    .A_7       (addKernel_36_A_7[31:0]), //i
    .A_8       (addKernel_36_A_8[31:0]), //i
    .S         (addKernel_36_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_37 (
    .A_0       (addKernel_37_A_0[31:0]), //i
    .A_1       (addKernel_37_A_1[31:0]), //i
    .A_2       (addKernel_37_A_2[31:0]), //i
    .A_3       (addKernel_37_A_3[31:0]), //i
    .A_4       (addKernel_37_A_4[31:0]), //i
    .A_5       (addKernel_37_A_5[31:0]), //i
    .A_6       (addKernel_37_A_6[31:0]), //i
    .A_7       (addKernel_37_A_7[31:0]), //i
    .A_8       (addKernel_37_A_8[31:0]), //i
    .S         (addKernel_37_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_38 (
    .A_0       (addKernel_38_A_0[31:0]), //i
    .A_1       (addKernel_38_A_1[31:0]), //i
    .A_2       (addKernel_38_A_2[31:0]), //i
    .A_3       (addKernel_38_A_3[31:0]), //i
    .A_4       (addKernel_38_A_4[31:0]), //i
    .A_5       (addKernel_38_A_5[31:0]), //i
    .A_6       (addKernel_38_A_6[31:0]), //i
    .A_7       (addKernel_38_A_7[31:0]), //i
    .A_8       (addKernel_38_A_8[31:0]), //i
    .S         (addKernel_38_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_39 (
    .A_0       (addKernel_39_A_0[31:0]), //i
    .A_1       (addKernel_39_A_1[31:0]), //i
    .A_2       (addKernel_39_A_2[31:0]), //i
    .A_3       (addKernel_39_A_3[31:0]), //i
    .A_4       (addKernel_39_A_4[31:0]), //i
    .A_5       (addKernel_39_A_5[31:0]), //i
    .A_6       (addKernel_39_A_6[31:0]), //i
    .A_7       (addKernel_39_A_7[31:0]), //i
    .A_8       (addKernel_39_A_8[31:0]), //i
    .S         (addKernel_39_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_40 (
    .A_0       (addKernel_40_A_0[31:0]), //i
    .A_1       (addKernel_40_A_1[31:0]), //i
    .A_2       (addKernel_40_A_2[31:0]), //i
    .A_3       (addKernel_40_A_3[31:0]), //i
    .A_4       (addKernel_40_A_4[31:0]), //i
    .A_5       (addKernel_40_A_5[31:0]), //i
    .A_6       (addKernel_40_A_6[31:0]), //i
    .A_7       (addKernel_40_A_7[31:0]), //i
    .A_8       (addKernel_40_A_8[31:0]), //i
    .S         (addKernel_40_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_41 (
    .A_0       (addKernel_41_A_0[31:0]), //i
    .A_1       (addKernel_41_A_1[31:0]), //i
    .A_2       (addKernel_41_A_2[31:0]), //i
    .A_3       (addKernel_41_A_3[31:0]), //i
    .A_4       (addKernel_41_A_4[31:0]), //i
    .A_5       (addKernel_41_A_5[31:0]), //i
    .A_6       (addKernel_41_A_6[31:0]), //i
    .A_7       (addKernel_41_A_7[31:0]), //i
    .A_8       (addKernel_41_A_8[31:0]), //i
    .S         (addKernel_41_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_42 (
    .A_0       (addKernel_42_A_0[31:0]), //i
    .A_1       (addKernel_42_A_1[31:0]), //i
    .A_2       (addKernel_42_A_2[31:0]), //i
    .A_3       (addKernel_42_A_3[31:0]), //i
    .A_4       (addKernel_42_A_4[31:0]), //i
    .A_5       (addKernel_42_A_5[31:0]), //i
    .A_6       (addKernel_42_A_6[31:0]), //i
    .A_7       (addKernel_42_A_7[31:0]), //i
    .A_8       (addKernel_42_A_8[31:0]), //i
    .S         (addKernel_42_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_43 (
    .A_0       (addKernel_43_A_0[31:0]), //i
    .A_1       (addKernel_43_A_1[31:0]), //i
    .A_2       (addKernel_43_A_2[31:0]), //i
    .A_3       (addKernel_43_A_3[31:0]), //i
    .A_4       (addKernel_43_A_4[31:0]), //i
    .A_5       (addKernel_43_A_5[31:0]), //i
    .A_6       (addKernel_43_A_6[31:0]), //i
    .A_7       (addKernel_43_A_7[31:0]), //i
    .A_8       (addKernel_43_A_8[31:0]), //i
    .S         (addKernel_43_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_44 (
    .A_0       (addKernel_44_A_0[31:0]), //i
    .A_1       (addKernel_44_A_1[31:0]), //i
    .A_2       (addKernel_44_A_2[31:0]), //i
    .A_3       (addKernel_44_A_3[31:0]), //i
    .A_4       (addKernel_44_A_4[31:0]), //i
    .A_5       (addKernel_44_A_5[31:0]), //i
    .A_6       (addKernel_44_A_6[31:0]), //i
    .A_7       (addKernel_44_A_7[31:0]), //i
    .A_8       (addKernel_44_A_8[31:0]), //i
    .S         (addKernel_44_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_45 (
    .A_0       (addKernel_45_A_0[31:0]), //i
    .A_1       (addKernel_45_A_1[31:0]), //i
    .A_2       (addKernel_45_A_2[31:0]), //i
    .A_3       (addKernel_45_A_3[31:0]), //i
    .A_4       (addKernel_45_A_4[31:0]), //i
    .A_5       (addKernel_45_A_5[31:0]), //i
    .A_6       (addKernel_45_A_6[31:0]), //i
    .A_7       (addKernel_45_A_7[31:0]), //i
    .A_8       (addKernel_45_A_8[31:0]), //i
    .S         (addKernel_45_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_46 (
    .A_0       (addKernel_46_A_0[31:0]), //i
    .A_1       (addKernel_46_A_1[31:0]), //i
    .A_2       (addKernel_46_A_2[31:0]), //i
    .A_3       (addKernel_46_A_3[31:0]), //i
    .A_4       (addKernel_46_A_4[31:0]), //i
    .A_5       (addKernel_46_A_5[31:0]), //i
    .A_6       (addKernel_46_A_6[31:0]), //i
    .A_7       (addKernel_46_A_7[31:0]), //i
    .A_8       (addKernel_46_A_8[31:0]), //i
    .S         (addKernel_46_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_47 (
    .A_0       (addKernel_47_A_0[31:0]), //i
    .A_1       (addKernel_47_A_1[31:0]), //i
    .A_2       (addKernel_47_A_2[31:0]), //i
    .A_3       (addKernel_47_A_3[31:0]), //i
    .A_4       (addKernel_47_A_4[31:0]), //i
    .A_5       (addKernel_47_A_5[31:0]), //i
    .A_6       (addKernel_47_A_6[31:0]), //i
    .A_7       (addKernel_47_A_7[31:0]), //i
    .A_8       (addKernel_47_A_8[31:0]), //i
    .S         (addKernel_47_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_48 (
    .A_0       (addKernel_48_A_0[31:0]), //i
    .A_1       (addKernel_48_A_1[31:0]), //i
    .A_2       (addKernel_48_A_2[31:0]), //i
    .A_3       (addKernel_48_A_3[31:0]), //i
    .A_4       (addKernel_48_A_4[31:0]), //i
    .A_5       (addKernel_48_A_5[31:0]), //i
    .A_6       (addKernel_48_A_6[31:0]), //i
    .A_7       (addKernel_48_A_7[31:0]), //i
    .A_8       (addKernel_48_A_8[31:0]), //i
    .S         (addKernel_48_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_49 (
    .A_0       (addKernel_49_A_0[31:0]), //i
    .A_1       (addKernel_49_A_1[31:0]), //i
    .A_2       (addKernel_49_A_2[31:0]), //i
    .A_3       (addKernel_49_A_3[31:0]), //i
    .A_4       (addKernel_49_A_4[31:0]), //i
    .A_5       (addKernel_49_A_5[31:0]), //i
    .A_6       (addKernel_49_A_6[31:0]), //i
    .A_7       (addKernel_49_A_7[31:0]), //i
    .A_8       (addKernel_49_A_8[31:0]), //i
    .S         (addKernel_49_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_50 (
    .A_0       (addKernel_50_A_0[31:0]), //i
    .A_1       (addKernel_50_A_1[31:0]), //i
    .A_2       (addKernel_50_A_2[31:0]), //i
    .A_3       (addKernel_50_A_3[31:0]), //i
    .A_4       (addKernel_50_A_4[31:0]), //i
    .A_5       (addKernel_50_A_5[31:0]), //i
    .A_6       (addKernel_50_A_6[31:0]), //i
    .A_7       (addKernel_50_A_7[31:0]), //i
    .A_8       (addKernel_50_A_8[31:0]), //i
    .S         (addKernel_50_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_51 (
    .A_0       (addKernel_51_A_0[31:0]), //i
    .A_1       (addKernel_51_A_1[31:0]), //i
    .A_2       (addKernel_51_A_2[31:0]), //i
    .A_3       (addKernel_51_A_3[31:0]), //i
    .A_4       (addKernel_51_A_4[31:0]), //i
    .A_5       (addKernel_51_A_5[31:0]), //i
    .A_6       (addKernel_51_A_6[31:0]), //i
    .A_7       (addKernel_51_A_7[31:0]), //i
    .A_8       (addKernel_51_A_8[31:0]), //i
    .S         (addKernel_51_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_52 (
    .A_0       (addKernel_52_A_0[31:0]), //i
    .A_1       (addKernel_52_A_1[31:0]), //i
    .A_2       (addKernel_52_A_2[31:0]), //i
    .A_3       (addKernel_52_A_3[31:0]), //i
    .A_4       (addKernel_52_A_4[31:0]), //i
    .A_5       (addKernel_52_A_5[31:0]), //i
    .A_6       (addKernel_52_A_6[31:0]), //i
    .A_7       (addKernel_52_A_7[31:0]), //i
    .A_8       (addKernel_52_A_8[31:0]), //i
    .S         (addKernel_52_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_53 (
    .A_0       (addKernel_53_A_0[31:0]), //i
    .A_1       (addKernel_53_A_1[31:0]), //i
    .A_2       (addKernel_53_A_2[31:0]), //i
    .A_3       (addKernel_53_A_3[31:0]), //i
    .A_4       (addKernel_53_A_4[31:0]), //i
    .A_5       (addKernel_53_A_5[31:0]), //i
    .A_6       (addKernel_53_A_6[31:0]), //i
    .A_7       (addKernel_53_A_7[31:0]), //i
    .A_8       (addKernel_53_A_8[31:0]), //i
    .S         (addKernel_53_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_54 (
    .A_0       (addKernel_54_A_0[31:0]), //i
    .A_1       (addKernel_54_A_1[31:0]), //i
    .A_2       (addKernel_54_A_2[31:0]), //i
    .A_3       (addKernel_54_A_3[31:0]), //i
    .A_4       (addKernel_54_A_4[31:0]), //i
    .A_5       (addKernel_54_A_5[31:0]), //i
    .A_6       (addKernel_54_A_6[31:0]), //i
    .A_7       (addKernel_54_A_7[31:0]), //i
    .A_8       (addKernel_54_A_8[31:0]), //i
    .S         (addKernel_54_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_55 (
    .A_0       (addKernel_55_A_0[31:0]), //i
    .A_1       (addKernel_55_A_1[31:0]), //i
    .A_2       (addKernel_55_A_2[31:0]), //i
    .A_3       (addKernel_55_A_3[31:0]), //i
    .A_4       (addKernel_55_A_4[31:0]), //i
    .A_5       (addKernel_55_A_5[31:0]), //i
    .A_6       (addKernel_55_A_6[31:0]), //i
    .A_7       (addKernel_55_A_7[31:0]), //i
    .A_8       (addKernel_55_A_8[31:0]), //i
    .S         (addKernel_55_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_56 (
    .A_0       (addKernel_56_A_0[31:0]), //i
    .A_1       (addKernel_56_A_1[31:0]), //i
    .A_2       (addKernel_56_A_2[31:0]), //i
    .A_3       (addKernel_56_A_3[31:0]), //i
    .A_4       (addKernel_56_A_4[31:0]), //i
    .A_5       (addKernel_56_A_5[31:0]), //i
    .A_6       (addKernel_56_A_6[31:0]), //i
    .A_7       (addKernel_56_A_7[31:0]), //i
    .A_8       (addKernel_56_A_8[31:0]), //i
    .S         (addKernel_56_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_57 (
    .A_0       (addKernel_57_A_0[31:0]), //i
    .A_1       (addKernel_57_A_1[31:0]), //i
    .A_2       (addKernel_57_A_2[31:0]), //i
    .A_3       (addKernel_57_A_3[31:0]), //i
    .A_4       (addKernel_57_A_4[31:0]), //i
    .A_5       (addKernel_57_A_5[31:0]), //i
    .A_6       (addKernel_57_A_6[31:0]), //i
    .A_7       (addKernel_57_A_7[31:0]), //i
    .A_8       (addKernel_57_A_8[31:0]), //i
    .S         (addKernel_57_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_58 (
    .A_0       (addKernel_58_A_0[31:0]), //i
    .A_1       (addKernel_58_A_1[31:0]), //i
    .A_2       (addKernel_58_A_2[31:0]), //i
    .A_3       (addKernel_58_A_3[31:0]), //i
    .A_4       (addKernel_58_A_4[31:0]), //i
    .A_5       (addKernel_58_A_5[31:0]), //i
    .A_6       (addKernel_58_A_6[31:0]), //i
    .A_7       (addKernel_58_A_7[31:0]), //i
    .A_8       (addKernel_58_A_8[31:0]), //i
    .S         (addKernel_58_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_59 (
    .A_0       (addKernel_59_A_0[31:0]), //i
    .A_1       (addKernel_59_A_1[31:0]), //i
    .A_2       (addKernel_59_A_2[31:0]), //i
    .A_3       (addKernel_59_A_3[31:0]), //i
    .A_4       (addKernel_59_A_4[31:0]), //i
    .A_5       (addKernel_59_A_5[31:0]), //i
    .A_6       (addKernel_59_A_6[31:0]), //i
    .A_7       (addKernel_59_A_7[31:0]), //i
    .A_8       (addKernel_59_A_8[31:0]), //i
    .S         (addKernel_59_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_60 (
    .A_0       (addKernel_60_A_0[31:0]), //i
    .A_1       (addKernel_60_A_1[31:0]), //i
    .A_2       (addKernel_60_A_2[31:0]), //i
    .A_3       (addKernel_60_A_3[31:0]), //i
    .A_4       (addKernel_60_A_4[31:0]), //i
    .A_5       (addKernel_60_A_5[31:0]), //i
    .A_6       (addKernel_60_A_6[31:0]), //i
    .A_7       (addKernel_60_A_7[31:0]), //i
    .A_8       (addKernel_60_A_8[31:0]), //i
    .S         (addKernel_60_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_61 (
    .A_0       (addKernel_61_A_0[31:0]), //i
    .A_1       (addKernel_61_A_1[31:0]), //i
    .A_2       (addKernel_61_A_2[31:0]), //i
    .A_3       (addKernel_61_A_3[31:0]), //i
    .A_4       (addKernel_61_A_4[31:0]), //i
    .A_5       (addKernel_61_A_5[31:0]), //i
    .A_6       (addKernel_61_A_6[31:0]), //i
    .A_7       (addKernel_61_A_7[31:0]), //i
    .A_8       (addKernel_61_A_8[31:0]), //i
    .S         (addKernel_61_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_62 (
    .A_0       (addKernel_62_A_0[31:0]), //i
    .A_1       (addKernel_62_A_1[31:0]), //i
    .A_2       (addKernel_62_A_2[31:0]), //i
    .A_3       (addKernel_62_A_3[31:0]), //i
    .A_4       (addKernel_62_A_4[31:0]), //i
    .A_5       (addKernel_62_A_5[31:0]), //i
    .A_6       (addKernel_62_A_6[31:0]), //i
    .A_7       (addKernel_62_A_7[31:0]), //i
    .A_8       (addKernel_62_A_8[31:0]), //i
    .S         (addKernel_62_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_63 (
    .A_0       (addKernel_63_A_0[31:0]), //i
    .A_1       (addKernel_63_A_1[31:0]), //i
    .A_2       (addKernel_63_A_2[31:0]), //i
    .A_3       (addKernel_63_A_3[31:0]), //i
    .A_4       (addKernel_63_A_4[31:0]), //i
    .A_5       (addKernel_63_A_5[31:0]), //i
    .A_6       (addKernel_63_A_6[31:0]), //i
    .A_7       (addKernel_63_A_7[31:0]), //i
    .A_8       (addKernel_63_A_8[31:0]), //i
    .S         (addKernel_63_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_64 (
    .A_0       (addKernel_64_A_0[31:0]), //i
    .A_1       (addKernel_64_A_1[31:0]), //i
    .A_2       (addKernel_64_A_2[31:0]), //i
    .A_3       (addKernel_64_A_3[31:0]), //i
    .A_4       (addKernel_64_A_4[31:0]), //i
    .A_5       (addKernel_64_A_5[31:0]), //i
    .A_6       (addKernel_64_A_6[31:0]), //i
    .A_7       (addKernel_64_A_7[31:0]), //i
    .A_8       (addKernel_64_A_8[31:0]), //i
    .S         (addKernel_64_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_65 (
    .A_0       (addKernel_65_A_0[31:0]), //i
    .A_1       (addKernel_65_A_1[31:0]), //i
    .A_2       (addKernel_65_A_2[31:0]), //i
    .A_3       (addKernel_65_A_3[31:0]), //i
    .A_4       (addKernel_65_A_4[31:0]), //i
    .A_5       (addKernel_65_A_5[31:0]), //i
    .A_6       (addKernel_65_A_6[31:0]), //i
    .A_7       (addKernel_65_A_7[31:0]), //i
    .A_8       (addKernel_65_A_8[31:0]), //i
    .S         (addKernel_65_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_66 (
    .A_0       (addKernel_66_A_0[31:0]), //i
    .A_1       (addKernel_66_A_1[31:0]), //i
    .A_2       (addKernel_66_A_2[31:0]), //i
    .A_3       (addKernel_66_A_3[31:0]), //i
    .A_4       (addKernel_66_A_4[31:0]), //i
    .A_5       (addKernel_66_A_5[31:0]), //i
    .A_6       (addKernel_66_A_6[31:0]), //i
    .A_7       (addKernel_66_A_7[31:0]), //i
    .A_8       (addKernel_66_A_8[31:0]), //i
    .S         (addKernel_66_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_67 (
    .A_0       (addKernel_67_A_0[31:0]), //i
    .A_1       (addKernel_67_A_1[31:0]), //i
    .A_2       (addKernel_67_A_2[31:0]), //i
    .A_3       (addKernel_67_A_3[31:0]), //i
    .A_4       (addKernel_67_A_4[31:0]), //i
    .A_5       (addKernel_67_A_5[31:0]), //i
    .A_6       (addKernel_67_A_6[31:0]), //i
    .A_7       (addKernel_67_A_7[31:0]), //i
    .A_8       (addKernel_67_A_8[31:0]), //i
    .S         (addKernel_67_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_68 (
    .A_0       (addKernel_68_A_0[31:0]), //i
    .A_1       (addKernel_68_A_1[31:0]), //i
    .A_2       (addKernel_68_A_2[31:0]), //i
    .A_3       (addKernel_68_A_3[31:0]), //i
    .A_4       (addKernel_68_A_4[31:0]), //i
    .A_5       (addKernel_68_A_5[31:0]), //i
    .A_6       (addKernel_68_A_6[31:0]), //i
    .A_7       (addKernel_68_A_7[31:0]), //i
    .A_8       (addKernel_68_A_8[31:0]), //i
    .S         (addKernel_68_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_69 (
    .A_0       (addKernel_69_A_0[31:0]), //i
    .A_1       (addKernel_69_A_1[31:0]), //i
    .A_2       (addKernel_69_A_2[31:0]), //i
    .A_3       (addKernel_69_A_3[31:0]), //i
    .A_4       (addKernel_69_A_4[31:0]), //i
    .A_5       (addKernel_69_A_5[31:0]), //i
    .A_6       (addKernel_69_A_6[31:0]), //i
    .A_7       (addKernel_69_A_7[31:0]), //i
    .A_8       (addKernel_69_A_8[31:0]), //i
    .S         (addKernel_69_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_70 (
    .A_0       (addKernel_70_A_0[31:0]), //i
    .A_1       (addKernel_70_A_1[31:0]), //i
    .A_2       (addKernel_70_A_2[31:0]), //i
    .A_3       (addKernel_70_A_3[31:0]), //i
    .A_4       (addKernel_70_A_4[31:0]), //i
    .A_5       (addKernel_70_A_5[31:0]), //i
    .A_6       (addKernel_70_A_6[31:0]), //i
    .A_7       (addKernel_70_A_7[31:0]), //i
    .A_8       (addKernel_70_A_8[31:0]), //i
    .S         (addKernel_70_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_71 (
    .A_0       (addKernel_71_A_0[31:0]), //i
    .A_1       (addKernel_71_A_1[31:0]), //i
    .A_2       (addKernel_71_A_2[31:0]), //i
    .A_3       (addKernel_71_A_3[31:0]), //i
    .A_4       (addKernel_71_A_4[31:0]), //i
    .A_5       (addKernel_71_A_5[31:0]), //i
    .A_6       (addKernel_71_A_6[31:0]), //i
    .A_7       (addKernel_71_A_7[31:0]), //i
    .A_8       (addKernel_71_A_8[31:0]), //i
    .S         (addKernel_71_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_72 (
    .A_0       (addKernel_72_A_0[31:0]), //i
    .A_1       (addKernel_72_A_1[31:0]), //i
    .A_2       (addKernel_72_A_2[31:0]), //i
    .A_3       (addKernel_72_A_3[31:0]), //i
    .A_4       (addKernel_72_A_4[31:0]), //i
    .A_5       (addKernel_72_A_5[31:0]), //i
    .A_6       (addKernel_72_A_6[31:0]), //i
    .A_7       (addKernel_72_A_7[31:0]), //i
    .A_8       (addKernel_72_A_8[31:0]), //i
    .S         (addKernel_72_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_73 (
    .A_0       (addKernel_73_A_0[31:0]), //i
    .A_1       (addKernel_73_A_1[31:0]), //i
    .A_2       (addKernel_73_A_2[31:0]), //i
    .A_3       (addKernel_73_A_3[31:0]), //i
    .A_4       (addKernel_73_A_4[31:0]), //i
    .A_5       (addKernel_73_A_5[31:0]), //i
    .A_6       (addKernel_73_A_6[31:0]), //i
    .A_7       (addKernel_73_A_7[31:0]), //i
    .A_8       (addKernel_73_A_8[31:0]), //i
    .S         (addKernel_73_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_74 (
    .A_0       (addKernel_74_A_0[31:0]), //i
    .A_1       (addKernel_74_A_1[31:0]), //i
    .A_2       (addKernel_74_A_2[31:0]), //i
    .A_3       (addKernel_74_A_3[31:0]), //i
    .A_4       (addKernel_74_A_4[31:0]), //i
    .A_5       (addKernel_74_A_5[31:0]), //i
    .A_6       (addKernel_74_A_6[31:0]), //i
    .A_7       (addKernel_74_A_7[31:0]), //i
    .A_8       (addKernel_74_A_8[31:0]), //i
    .S         (addKernel_74_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_75 (
    .A_0       (addKernel_75_A_0[31:0]), //i
    .A_1       (addKernel_75_A_1[31:0]), //i
    .A_2       (addKernel_75_A_2[31:0]), //i
    .A_3       (addKernel_75_A_3[31:0]), //i
    .A_4       (addKernel_75_A_4[31:0]), //i
    .A_5       (addKernel_75_A_5[31:0]), //i
    .A_6       (addKernel_75_A_6[31:0]), //i
    .A_7       (addKernel_75_A_7[31:0]), //i
    .A_8       (addKernel_75_A_8[31:0]), //i
    .S         (addKernel_75_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_76 (
    .A_0       (addKernel_76_A_0[31:0]), //i
    .A_1       (addKernel_76_A_1[31:0]), //i
    .A_2       (addKernel_76_A_2[31:0]), //i
    .A_3       (addKernel_76_A_3[31:0]), //i
    .A_4       (addKernel_76_A_4[31:0]), //i
    .A_5       (addKernel_76_A_5[31:0]), //i
    .A_6       (addKernel_76_A_6[31:0]), //i
    .A_7       (addKernel_76_A_7[31:0]), //i
    .A_8       (addKernel_76_A_8[31:0]), //i
    .S         (addKernel_76_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_77 (
    .A_0       (addKernel_77_A_0[31:0]), //i
    .A_1       (addKernel_77_A_1[31:0]), //i
    .A_2       (addKernel_77_A_2[31:0]), //i
    .A_3       (addKernel_77_A_3[31:0]), //i
    .A_4       (addKernel_77_A_4[31:0]), //i
    .A_5       (addKernel_77_A_5[31:0]), //i
    .A_6       (addKernel_77_A_6[31:0]), //i
    .A_7       (addKernel_77_A_7[31:0]), //i
    .A_8       (addKernel_77_A_8[31:0]), //i
    .S         (addKernel_77_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_78 (
    .A_0       (addKernel_78_A_0[31:0]), //i
    .A_1       (addKernel_78_A_1[31:0]), //i
    .A_2       (addKernel_78_A_2[31:0]), //i
    .A_3       (addKernel_78_A_3[31:0]), //i
    .A_4       (addKernel_78_A_4[31:0]), //i
    .A_5       (addKernel_78_A_5[31:0]), //i
    .A_6       (addKernel_78_A_6[31:0]), //i
    .A_7       (addKernel_78_A_7[31:0]), //i
    .A_8       (addKernel_78_A_8[31:0]), //i
    .S         (addKernel_78_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_79 (
    .A_0       (addKernel_79_A_0[31:0]), //i
    .A_1       (addKernel_79_A_1[31:0]), //i
    .A_2       (addKernel_79_A_2[31:0]), //i
    .A_3       (addKernel_79_A_3[31:0]), //i
    .A_4       (addKernel_79_A_4[31:0]), //i
    .A_5       (addKernel_79_A_5[31:0]), //i
    .A_6       (addKernel_79_A_6[31:0]), //i
    .A_7       (addKernel_79_A_7[31:0]), //i
    .A_8       (addKernel_79_A_8[31:0]), //i
    .S         (addKernel_79_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_80 (
    .A_0       (addKernel_80_A_0[31:0]), //i
    .A_1       (addKernel_80_A_1[31:0]), //i
    .A_2       (addKernel_80_A_2[31:0]), //i
    .A_3       (addKernel_80_A_3[31:0]), //i
    .A_4       (addKernel_80_A_4[31:0]), //i
    .A_5       (addKernel_80_A_5[31:0]), //i
    .A_6       (addKernel_80_A_6[31:0]), //i
    .A_7       (addKernel_80_A_7[31:0]), //i
    .A_8       (addKernel_80_A_8[31:0]), //i
    .S         (addKernel_80_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_81 (
    .A_0       (addKernel_81_A_0[31:0]), //i
    .A_1       (addKernel_81_A_1[31:0]), //i
    .A_2       (addKernel_81_A_2[31:0]), //i
    .A_3       (addKernel_81_A_3[31:0]), //i
    .A_4       (addKernel_81_A_4[31:0]), //i
    .A_5       (addKernel_81_A_5[31:0]), //i
    .A_6       (addKernel_81_A_6[31:0]), //i
    .A_7       (addKernel_81_A_7[31:0]), //i
    .A_8       (addKernel_81_A_8[31:0]), //i
    .S         (addKernel_81_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_82 (
    .A_0       (addKernel_82_A_0[31:0]), //i
    .A_1       (addKernel_82_A_1[31:0]), //i
    .A_2       (addKernel_82_A_2[31:0]), //i
    .A_3       (addKernel_82_A_3[31:0]), //i
    .A_4       (addKernel_82_A_4[31:0]), //i
    .A_5       (addKernel_82_A_5[31:0]), //i
    .A_6       (addKernel_82_A_6[31:0]), //i
    .A_7       (addKernel_82_A_7[31:0]), //i
    .A_8       (addKernel_82_A_8[31:0]), //i
    .S         (addKernel_82_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_83 (
    .A_0       (addKernel_83_A_0[31:0]), //i
    .A_1       (addKernel_83_A_1[31:0]), //i
    .A_2       (addKernel_83_A_2[31:0]), //i
    .A_3       (addKernel_83_A_3[31:0]), //i
    .A_4       (addKernel_83_A_4[31:0]), //i
    .A_5       (addKernel_83_A_5[31:0]), //i
    .A_6       (addKernel_83_A_6[31:0]), //i
    .A_7       (addKernel_83_A_7[31:0]), //i
    .A_8       (addKernel_83_A_8[31:0]), //i
    .S         (addKernel_83_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_84 (
    .A_0       (addKernel_84_A_0[31:0]), //i
    .A_1       (addKernel_84_A_1[31:0]), //i
    .A_2       (addKernel_84_A_2[31:0]), //i
    .A_3       (addKernel_84_A_3[31:0]), //i
    .A_4       (addKernel_84_A_4[31:0]), //i
    .A_5       (addKernel_84_A_5[31:0]), //i
    .A_6       (addKernel_84_A_6[31:0]), //i
    .A_7       (addKernel_84_A_7[31:0]), //i
    .A_8       (addKernel_84_A_8[31:0]), //i
    .S         (addKernel_84_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_85 (
    .A_0       (addKernel_85_A_0[31:0]), //i
    .A_1       (addKernel_85_A_1[31:0]), //i
    .A_2       (addKernel_85_A_2[31:0]), //i
    .A_3       (addKernel_85_A_3[31:0]), //i
    .A_4       (addKernel_85_A_4[31:0]), //i
    .A_5       (addKernel_85_A_5[31:0]), //i
    .A_6       (addKernel_85_A_6[31:0]), //i
    .A_7       (addKernel_85_A_7[31:0]), //i
    .A_8       (addKernel_85_A_8[31:0]), //i
    .S         (addKernel_85_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_86 (
    .A_0       (addKernel_86_A_0[31:0]), //i
    .A_1       (addKernel_86_A_1[31:0]), //i
    .A_2       (addKernel_86_A_2[31:0]), //i
    .A_3       (addKernel_86_A_3[31:0]), //i
    .A_4       (addKernel_86_A_4[31:0]), //i
    .A_5       (addKernel_86_A_5[31:0]), //i
    .A_6       (addKernel_86_A_6[31:0]), //i
    .A_7       (addKernel_86_A_7[31:0]), //i
    .A_8       (addKernel_86_A_8[31:0]), //i
    .S         (addKernel_86_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_87 (
    .A_0       (addKernel_87_A_0[31:0]), //i
    .A_1       (addKernel_87_A_1[31:0]), //i
    .A_2       (addKernel_87_A_2[31:0]), //i
    .A_3       (addKernel_87_A_3[31:0]), //i
    .A_4       (addKernel_87_A_4[31:0]), //i
    .A_5       (addKernel_87_A_5[31:0]), //i
    .A_6       (addKernel_87_A_6[31:0]), //i
    .A_7       (addKernel_87_A_7[31:0]), //i
    .A_8       (addKernel_87_A_8[31:0]), //i
    .S         (addKernel_87_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_88 (
    .A_0       (addKernel_88_A_0[31:0]), //i
    .A_1       (addKernel_88_A_1[31:0]), //i
    .A_2       (addKernel_88_A_2[31:0]), //i
    .A_3       (addKernel_88_A_3[31:0]), //i
    .A_4       (addKernel_88_A_4[31:0]), //i
    .A_5       (addKernel_88_A_5[31:0]), //i
    .A_6       (addKernel_88_A_6[31:0]), //i
    .A_7       (addKernel_88_A_7[31:0]), //i
    .A_8       (addKernel_88_A_8[31:0]), //i
    .S         (addKernel_88_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_89 (
    .A_0       (addKernel_89_A_0[31:0]), //i
    .A_1       (addKernel_89_A_1[31:0]), //i
    .A_2       (addKernel_89_A_2[31:0]), //i
    .A_3       (addKernel_89_A_3[31:0]), //i
    .A_4       (addKernel_89_A_4[31:0]), //i
    .A_5       (addKernel_89_A_5[31:0]), //i
    .A_6       (addKernel_89_A_6[31:0]), //i
    .A_7       (addKernel_89_A_7[31:0]), //i
    .A_8       (addKernel_89_A_8[31:0]), //i
    .S         (addKernel_89_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_90 (
    .A_0       (addKernel_90_A_0[31:0]), //i
    .A_1       (addKernel_90_A_1[31:0]), //i
    .A_2       (addKernel_90_A_2[31:0]), //i
    .A_3       (addKernel_90_A_3[31:0]), //i
    .A_4       (addKernel_90_A_4[31:0]), //i
    .A_5       (addKernel_90_A_5[31:0]), //i
    .A_6       (addKernel_90_A_6[31:0]), //i
    .A_7       (addKernel_90_A_7[31:0]), //i
    .A_8       (addKernel_90_A_8[31:0]), //i
    .S         (addKernel_90_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_91 (
    .A_0       (addKernel_91_A_0[31:0]), //i
    .A_1       (addKernel_91_A_1[31:0]), //i
    .A_2       (addKernel_91_A_2[31:0]), //i
    .A_3       (addKernel_91_A_3[31:0]), //i
    .A_4       (addKernel_91_A_4[31:0]), //i
    .A_5       (addKernel_91_A_5[31:0]), //i
    .A_6       (addKernel_91_A_6[31:0]), //i
    .A_7       (addKernel_91_A_7[31:0]), //i
    .A_8       (addKernel_91_A_8[31:0]), //i
    .S         (addKernel_91_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_92 (
    .A_0       (addKernel_92_A_0[31:0]), //i
    .A_1       (addKernel_92_A_1[31:0]), //i
    .A_2       (addKernel_92_A_2[31:0]), //i
    .A_3       (addKernel_92_A_3[31:0]), //i
    .A_4       (addKernel_92_A_4[31:0]), //i
    .A_5       (addKernel_92_A_5[31:0]), //i
    .A_6       (addKernel_92_A_6[31:0]), //i
    .A_7       (addKernel_92_A_7[31:0]), //i
    .A_8       (addKernel_92_A_8[31:0]), //i
    .S         (addKernel_92_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_93 (
    .A_0       (addKernel_93_A_0[31:0]), //i
    .A_1       (addKernel_93_A_1[31:0]), //i
    .A_2       (addKernel_93_A_2[31:0]), //i
    .A_3       (addKernel_93_A_3[31:0]), //i
    .A_4       (addKernel_93_A_4[31:0]), //i
    .A_5       (addKernel_93_A_5[31:0]), //i
    .A_6       (addKernel_93_A_6[31:0]), //i
    .A_7       (addKernel_93_A_7[31:0]), //i
    .A_8       (addKernel_93_A_8[31:0]), //i
    .S         (addKernel_93_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_94 (
    .A_0       (addKernel_94_A_0[31:0]), //i
    .A_1       (addKernel_94_A_1[31:0]), //i
    .A_2       (addKernel_94_A_2[31:0]), //i
    .A_3       (addKernel_94_A_3[31:0]), //i
    .A_4       (addKernel_94_A_4[31:0]), //i
    .A_5       (addKernel_94_A_5[31:0]), //i
    .A_6       (addKernel_94_A_6[31:0]), //i
    .A_7       (addKernel_94_A_7[31:0]), //i
    .A_8       (addKernel_94_A_8[31:0]), //i
    .S         (addKernel_94_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_95 (
    .A_0       (addKernel_95_A_0[31:0]), //i
    .A_1       (addKernel_95_A_1[31:0]), //i
    .A_2       (addKernel_95_A_2[31:0]), //i
    .A_3       (addKernel_95_A_3[31:0]), //i
    .A_4       (addKernel_95_A_4[31:0]), //i
    .A_5       (addKernel_95_A_5[31:0]), //i
    .A_6       (addKernel_95_A_6[31:0]), //i
    .A_7       (addKernel_95_A_7[31:0]), //i
    .A_8       (addKernel_95_A_8[31:0]), //i
    .S         (addKernel_95_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_96 (
    .A_0       (addKernel_96_A_0[31:0]), //i
    .A_1       (addKernel_96_A_1[31:0]), //i
    .A_2       (addKernel_96_A_2[31:0]), //i
    .A_3       (addKernel_96_A_3[31:0]), //i
    .A_4       (addKernel_96_A_4[31:0]), //i
    .A_5       (addKernel_96_A_5[31:0]), //i
    .A_6       (addKernel_96_A_6[31:0]), //i
    .A_7       (addKernel_96_A_7[31:0]), //i
    .A_8       (addKernel_96_A_8[31:0]), //i
    .S         (addKernel_96_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_97 (
    .A_0       (addKernel_97_A_0[31:0]), //i
    .A_1       (addKernel_97_A_1[31:0]), //i
    .A_2       (addKernel_97_A_2[31:0]), //i
    .A_3       (addKernel_97_A_3[31:0]), //i
    .A_4       (addKernel_97_A_4[31:0]), //i
    .A_5       (addKernel_97_A_5[31:0]), //i
    .A_6       (addKernel_97_A_6[31:0]), //i
    .A_7       (addKernel_97_A_7[31:0]), //i
    .A_8       (addKernel_97_A_8[31:0]), //i
    .S         (addKernel_97_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_98 (
    .A_0       (addKernel_98_A_0[31:0]), //i
    .A_1       (addKernel_98_A_1[31:0]), //i
    .A_2       (addKernel_98_A_2[31:0]), //i
    .A_3       (addKernel_98_A_3[31:0]), //i
    .A_4       (addKernel_98_A_4[31:0]), //i
    .A_5       (addKernel_98_A_5[31:0]), //i
    .A_6       (addKernel_98_A_6[31:0]), //i
    .A_7       (addKernel_98_A_7[31:0]), //i
    .A_8       (addKernel_98_A_8[31:0]), //i
    .S         (addKernel_98_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_99 (
    .A_0       (addKernel_99_A_0[31:0]), //i
    .A_1       (addKernel_99_A_1[31:0]), //i
    .A_2       (addKernel_99_A_2[31:0]), //i
    .A_3       (addKernel_99_A_3[31:0]), //i
    .A_4       (addKernel_99_A_4[31:0]), //i
    .A_5       (addKernel_99_A_5[31:0]), //i
    .A_6       (addKernel_99_A_6[31:0]), //i
    .A_7       (addKernel_99_A_7[31:0]), //i
    .A_8       (addKernel_99_A_8[31:0]), //i
    .S         (addKernel_99_S[39:0]  ), //o
    .clk       (clk                   ), //i
    .reset     (reset                 ), //i
    .softReset (softReset             )  //i
  );
  xAddTimes addKernel_100 (
    .A_0       (addKernel_100_A_0[31:0]), //i
    .A_1       (addKernel_100_A_1[31:0]), //i
    .A_2       (addKernel_100_A_2[31:0]), //i
    .A_3       (addKernel_100_A_3[31:0]), //i
    .A_4       (addKernel_100_A_4[31:0]), //i
    .A_5       (addKernel_100_A_5[31:0]), //i
    .A_6       (addKernel_100_A_6[31:0]), //i
    .A_7       (addKernel_100_A_7[31:0]), //i
    .A_8       (addKernel_100_A_8[31:0]), //i
    .S         (addKernel_100_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_101 (
    .A_0       (addKernel_101_A_0[31:0]), //i
    .A_1       (addKernel_101_A_1[31:0]), //i
    .A_2       (addKernel_101_A_2[31:0]), //i
    .A_3       (addKernel_101_A_3[31:0]), //i
    .A_4       (addKernel_101_A_4[31:0]), //i
    .A_5       (addKernel_101_A_5[31:0]), //i
    .A_6       (addKernel_101_A_6[31:0]), //i
    .A_7       (addKernel_101_A_7[31:0]), //i
    .A_8       (addKernel_101_A_8[31:0]), //i
    .S         (addKernel_101_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_102 (
    .A_0       (addKernel_102_A_0[31:0]), //i
    .A_1       (addKernel_102_A_1[31:0]), //i
    .A_2       (addKernel_102_A_2[31:0]), //i
    .A_3       (addKernel_102_A_3[31:0]), //i
    .A_4       (addKernel_102_A_4[31:0]), //i
    .A_5       (addKernel_102_A_5[31:0]), //i
    .A_6       (addKernel_102_A_6[31:0]), //i
    .A_7       (addKernel_102_A_7[31:0]), //i
    .A_8       (addKernel_102_A_8[31:0]), //i
    .S         (addKernel_102_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_103 (
    .A_0       (addKernel_103_A_0[31:0]), //i
    .A_1       (addKernel_103_A_1[31:0]), //i
    .A_2       (addKernel_103_A_2[31:0]), //i
    .A_3       (addKernel_103_A_3[31:0]), //i
    .A_4       (addKernel_103_A_4[31:0]), //i
    .A_5       (addKernel_103_A_5[31:0]), //i
    .A_6       (addKernel_103_A_6[31:0]), //i
    .A_7       (addKernel_103_A_7[31:0]), //i
    .A_8       (addKernel_103_A_8[31:0]), //i
    .S         (addKernel_103_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_104 (
    .A_0       (addKernel_104_A_0[31:0]), //i
    .A_1       (addKernel_104_A_1[31:0]), //i
    .A_2       (addKernel_104_A_2[31:0]), //i
    .A_3       (addKernel_104_A_3[31:0]), //i
    .A_4       (addKernel_104_A_4[31:0]), //i
    .A_5       (addKernel_104_A_5[31:0]), //i
    .A_6       (addKernel_104_A_6[31:0]), //i
    .A_7       (addKernel_104_A_7[31:0]), //i
    .A_8       (addKernel_104_A_8[31:0]), //i
    .S         (addKernel_104_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_105 (
    .A_0       (addKernel_105_A_0[31:0]), //i
    .A_1       (addKernel_105_A_1[31:0]), //i
    .A_2       (addKernel_105_A_2[31:0]), //i
    .A_3       (addKernel_105_A_3[31:0]), //i
    .A_4       (addKernel_105_A_4[31:0]), //i
    .A_5       (addKernel_105_A_5[31:0]), //i
    .A_6       (addKernel_105_A_6[31:0]), //i
    .A_7       (addKernel_105_A_7[31:0]), //i
    .A_8       (addKernel_105_A_8[31:0]), //i
    .S         (addKernel_105_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_106 (
    .A_0       (addKernel_106_A_0[31:0]), //i
    .A_1       (addKernel_106_A_1[31:0]), //i
    .A_2       (addKernel_106_A_2[31:0]), //i
    .A_3       (addKernel_106_A_3[31:0]), //i
    .A_4       (addKernel_106_A_4[31:0]), //i
    .A_5       (addKernel_106_A_5[31:0]), //i
    .A_6       (addKernel_106_A_6[31:0]), //i
    .A_7       (addKernel_106_A_7[31:0]), //i
    .A_8       (addKernel_106_A_8[31:0]), //i
    .S         (addKernel_106_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_107 (
    .A_0       (addKernel_107_A_0[31:0]), //i
    .A_1       (addKernel_107_A_1[31:0]), //i
    .A_2       (addKernel_107_A_2[31:0]), //i
    .A_3       (addKernel_107_A_3[31:0]), //i
    .A_4       (addKernel_107_A_4[31:0]), //i
    .A_5       (addKernel_107_A_5[31:0]), //i
    .A_6       (addKernel_107_A_6[31:0]), //i
    .A_7       (addKernel_107_A_7[31:0]), //i
    .A_8       (addKernel_107_A_8[31:0]), //i
    .S         (addKernel_107_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_108 (
    .A_0       (addKernel_108_A_0[31:0]), //i
    .A_1       (addKernel_108_A_1[31:0]), //i
    .A_2       (addKernel_108_A_2[31:0]), //i
    .A_3       (addKernel_108_A_3[31:0]), //i
    .A_4       (addKernel_108_A_4[31:0]), //i
    .A_5       (addKernel_108_A_5[31:0]), //i
    .A_6       (addKernel_108_A_6[31:0]), //i
    .A_7       (addKernel_108_A_7[31:0]), //i
    .A_8       (addKernel_108_A_8[31:0]), //i
    .S         (addKernel_108_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_109 (
    .A_0       (addKernel_109_A_0[31:0]), //i
    .A_1       (addKernel_109_A_1[31:0]), //i
    .A_2       (addKernel_109_A_2[31:0]), //i
    .A_3       (addKernel_109_A_3[31:0]), //i
    .A_4       (addKernel_109_A_4[31:0]), //i
    .A_5       (addKernel_109_A_5[31:0]), //i
    .A_6       (addKernel_109_A_6[31:0]), //i
    .A_7       (addKernel_109_A_7[31:0]), //i
    .A_8       (addKernel_109_A_8[31:0]), //i
    .S         (addKernel_109_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_110 (
    .A_0       (addKernel_110_A_0[31:0]), //i
    .A_1       (addKernel_110_A_1[31:0]), //i
    .A_2       (addKernel_110_A_2[31:0]), //i
    .A_3       (addKernel_110_A_3[31:0]), //i
    .A_4       (addKernel_110_A_4[31:0]), //i
    .A_5       (addKernel_110_A_5[31:0]), //i
    .A_6       (addKernel_110_A_6[31:0]), //i
    .A_7       (addKernel_110_A_7[31:0]), //i
    .A_8       (addKernel_110_A_8[31:0]), //i
    .S         (addKernel_110_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_111 (
    .A_0       (addKernel_111_A_0[31:0]), //i
    .A_1       (addKernel_111_A_1[31:0]), //i
    .A_2       (addKernel_111_A_2[31:0]), //i
    .A_3       (addKernel_111_A_3[31:0]), //i
    .A_4       (addKernel_111_A_4[31:0]), //i
    .A_5       (addKernel_111_A_5[31:0]), //i
    .A_6       (addKernel_111_A_6[31:0]), //i
    .A_7       (addKernel_111_A_7[31:0]), //i
    .A_8       (addKernel_111_A_8[31:0]), //i
    .S         (addKernel_111_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_112 (
    .A_0       (addKernel_112_A_0[31:0]), //i
    .A_1       (addKernel_112_A_1[31:0]), //i
    .A_2       (addKernel_112_A_2[31:0]), //i
    .A_3       (addKernel_112_A_3[31:0]), //i
    .A_4       (addKernel_112_A_4[31:0]), //i
    .A_5       (addKernel_112_A_5[31:0]), //i
    .A_6       (addKernel_112_A_6[31:0]), //i
    .A_7       (addKernel_112_A_7[31:0]), //i
    .A_8       (addKernel_112_A_8[31:0]), //i
    .S         (addKernel_112_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_113 (
    .A_0       (addKernel_113_A_0[31:0]), //i
    .A_1       (addKernel_113_A_1[31:0]), //i
    .A_2       (addKernel_113_A_2[31:0]), //i
    .A_3       (addKernel_113_A_3[31:0]), //i
    .A_4       (addKernel_113_A_4[31:0]), //i
    .A_5       (addKernel_113_A_5[31:0]), //i
    .A_6       (addKernel_113_A_6[31:0]), //i
    .A_7       (addKernel_113_A_7[31:0]), //i
    .A_8       (addKernel_113_A_8[31:0]), //i
    .S         (addKernel_113_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_114 (
    .A_0       (addKernel_114_A_0[31:0]), //i
    .A_1       (addKernel_114_A_1[31:0]), //i
    .A_2       (addKernel_114_A_2[31:0]), //i
    .A_3       (addKernel_114_A_3[31:0]), //i
    .A_4       (addKernel_114_A_4[31:0]), //i
    .A_5       (addKernel_114_A_5[31:0]), //i
    .A_6       (addKernel_114_A_6[31:0]), //i
    .A_7       (addKernel_114_A_7[31:0]), //i
    .A_8       (addKernel_114_A_8[31:0]), //i
    .S         (addKernel_114_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_115 (
    .A_0       (addKernel_115_A_0[31:0]), //i
    .A_1       (addKernel_115_A_1[31:0]), //i
    .A_2       (addKernel_115_A_2[31:0]), //i
    .A_3       (addKernel_115_A_3[31:0]), //i
    .A_4       (addKernel_115_A_4[31:0]), //i
    .A_5       (addKernel_115_A_5[31:0]), //i
    .A_6       (addKernel_115_A_6[31:0]), //i
    .A_7       (addKernel_115_A_7[31:0]), //i
    .A_8       (addKernel_115_A_8[31:0]), //i
    .S         (addKernel_115_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_116 (
    .A_0       (addKernel_116_A_0[31:0]), //i
    .A_1       (addKernel_116_A_1[31:0]), //i
    .A_2       (addKernel_116_A_2[31:0]), //i
    .A_3       (addKernel_116_A_3[31:0]), //i
    .A_4       (addKernel_116_A_4[31:0]), //i
    .A_5       (addKernel_116_A_5[31:0]), //i
    .A_6       (addKernel_116_A_6[31:0]), //i
    .A_7       (addKernel_116_A_7[31:0]), //i
    .A_8       (addKernel_116_A_8[31:0]), //i
    .S         (addKernel_116_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_117 (
    .A_0       (addKernel_117_A_0[31:0]), //i
    .A_1       (addKernel_117_A_1[31:0]), //i
    .A_2       (addKernel_117_A_2[31:0]), //i
    .A_3       (addKernel_117_A_3[31:0]), //i
    .A_4       (addKernel_117_A_4[31:0]), //i
    .A_5       (addKernel_117_A_5[31:0]), //i
    .A_6       (addKernel_117_A_6[31:0]), //i
    .A_7       (addKernel_117_A_7[31:0]), //i
    .A_8       (addKernel_117_A_8[31:0]), //i
    .S         (addKernel_117_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_118 (
    .A_0       (addKernel_118_A_0[31:0]), //i
    .A_1       (addKernel_118_A_1[31:0]), //i
    .A_2       (addKernel_118_A_2[31:0]), //i
    .A_3       (addKernel_118_A_3[31:0]), //i
    .A_4       (addKernel_118_A_4[31:0]), //i
    .A_5       (addKernel_118_A_5[31:0]), //i
    .A_6       (addKernel_118_A_6[31:0]), //i
    .A_7       (addKernel_118_A_7[31:0]), //i
    .A_8       (addKernel_118_A_8[31:0]), //i
    .S         (addKernel_118_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_119 (
    .A_0       (addKernel_119_A_0[31:0]), //i
    .A_1       (addKernel_119_A_1[31:0]), //i
    .A_2       (addKernel_119_A_2[31:0]), //i
    .A_3       (addKernel_119_A_3[31:0]), //i
    .A_4       (addKernel_119_A_4[31:0]), //i
    .A_5       (addKernel_119_A_5[31:0]), //i
    .A_6       (addKernel_119_A_6[31:0]), //i
    .A_7       (addKernel_119_A_7[31:0]), //i
    .A_8       (addKernel_119_A_8[31:0]), //i
    .S         (addKernel_119_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_120 (
    .A_0       (addKernel_120_A_0[31:0]), //i
    .A_1       (addKernel_120_A_1[31:0]), //i
    .A_2       (addKernel_120_A_2[31:0]), //i
    .A_3       (addKernel_120_A_3[31:0]), //i
    .A_4       (addKernel_120_A_4[31:0]), //i
    .A_5       (addKernel_120_A_5[31:0]), //i
    .A_6       (addKernel_120_A_6[31:0]), //i
    .A_7       (addKernel_120_A_7[31:0]), //i
    .A_8       (addKernel_120_A_8[31:0]), //i
    .S         (addKernel_120_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_121 (
    .A_0       (addKernel_121_A_0[31:0]), //i
    .A_1       (addKernel_121_A_1[31:0]), //i
    .A_2       (addKernel_121_A_2[31:0]), //i
    .A_3       (addKernel_121_A_3[31:0]), //i
    .A_4       (addKernel_121_A_4[31:0]), //i
    .A_5       (addKernel_121_A_5[31:0]), //i
    .A_6       (addKernel_121_A_6[31:0]), //i
    .A_7       (addKernel_121_A_7[31:0]), //i
    .A_8       (addKernel_121_A_8[31:0]), //i
    .S         (addKernel_121_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_122 (
    .A_0       (addKernel_122_A_0[31:0]), //i
    .A_1       (addKernel_122_A_1[31:0]), //i
    .A_2       (addKernel_122_A_2[31:0]), //i
    .A_3       (addKernel_122_A_3[31:0]), //i
    .A_4       (addKernel_122_A_4[31:0]), //i
    .A_5       (addKernel_122_A_5[31:0]), //i
    .A_6       (addKernel_122_A_6[31:0]), //i
    .A_7       (addKernel_122_A_7[31:0]), //i
    .A_8       (addKernel_122_A_8[31:0]), //i
    .S         (addKernel_122_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_123 (
    .A_0       (addKernel_123_A_0[31:0]), //i
    .A_1       (addKernel_123_A_1[31:0]), //i
    .A_2       (addKernel_123_A_2[31:0]), //i
    .A_3       (addKernel_123_A_3[31:0]), //i
    .A_4       (addKernel_123_A_4[31:0]), //i
    .A_5       (addKernel_123_A_5[31:0]), //i
    .A_6       (addKernel_123_A_6[31:0]), //i
    .A_7       (addKernel_123_A_7[31:0]), //i
    .A_8       (addKernel_123_A_8[31:0]), //i
    .S         (addKernel_123_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_124 (
    .A_0       (addKernel_124_A_0[31:0]), //i
    .A_1       (addKernel_124_A_1[31:0]), //i
    .A_2       (addKernel_124_A_2[31:0]), //i
    .A_3       (addKernel_124_A_3[31:0]), //i
    .A_4       (addKernel_124_A_4[31:0]), //i
    .A_5       (addKernel_124_A_5[31:0]), //i
    .A_6       (addKernel_124_A_6[31:0]), //i
    .A_7       (addKernel_124_A_7[31:0]), //i
    .A_8       (addKernel_124_A_8[31:0]), //i
    .S         (addKernel_124_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_125 (
    .A_0       (addKernel_125_A_0[31:0]), //i
    .A_1       (addKernel_125_A_1[31:0]), //i
    .A_2       (addKernel_125_A_2[31:0]), //i
    .A_3       (addKernel_125_A_3[31:0]), //i
    .A_4       (addKernel_125_A_4[31:0]), //i
    .A_5       (addKernel_125_A_5[31:0]), //i
    .A_6       (addKernel_125_A_6[31:0]), //i
    .A_7       (addKernel_125_A_7[31:0]), //i
    .A_8       (addKernel_125_A_8[31:0]), //i
    .S         (addKernel_125_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_126 (
    .A_0       (addKernel_126_A_0[31:0]), //i
    .A_1       (addKernel_126_A_1[31:0]), //i
    .A_2       (addKernel_126_A_2[31:0]), //i
    .A_3       (addKernel_126_A_3[31:0]), //i
    .A_4       (addKernel_126_A_4[31:0]), //i
    .A_5       (addKernel_126_A_5[31:0]), //i
    .A_6       (addKernel_126_A_6[31:0]), //i
    .A_7       (addKernel_126_A_7[31:0]), //i
    .A_8       (addKernel_126_A_8[31:0]), //i
    .S         (addKernel_126_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes addKernel_127 (
    .A_0       (addKernel_127_A_0[31:0]), //i
    .A_1       (addKernel_127_A_1[31:0]), //i
    .A_2       (addKernel_127_A_2[31:0]), //i
    .A_3       (addKernel_127_A_3[31:0]), //i
    .A_4       (addKernel_127_A_4[31:0]), //i
    .A_5       (addKernel_127_A_5[31:0]), //i
    .A_6       (addKernel_127_A_6[31:0]), //i
    .A_7       (addKernel_127_A_7[31:0]), //i
    .A_8       (addKernel_127_A_8[31:0]), //i
    .S         (addKernel_127_S[39:0]  ), //o
    .clk       (clk                    ), //i
    .reset     (reset                  ), //i
    .softReset (softReset              )  //i
  );
  xAddTimes_128 xAddTimes_136 (
    .A_0       (addKernel_S[39:0]    ), //i
    .A_1       (addKernel_1_S[39:0]  ), //i
    .A_2       (addKernel_2_S[39:0]  ), //i
    .A_3       (addKernel_3_S[39:0]  ), //i
    .A_4       (addKernel_4_S[39:0]  ), //i
    .A_5       (addKernel_5_S[39:0]  ), //i
    .A_6       (addKernel_6_S[39:0]  ), //i
    .A_7       (addKernel_7_S[39:0]  ), //i
    .A_8       (addKernel_8_S[39:0]  ), //i
    .A_9       (addKernel_9_S[39:0]  ), //i
    .A_10      (addKernel_10_S[39:0] ), //i
    .A_11      (addKernel_11_S[39:0] ), //i
    .A_12      (addKernel_12_S[39:0] ), //i
    .A_13      (addKernel_13_S[39:0] ), //i
    .A_14      (addKernel_14_S[39:0] ), //i
    .A_15      (addKernel_15_S[39:0] ), //i
    .S         (xAddTimes_136_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_137 (
    .A_0       (addKernel_16_S[39:0] ), //i
    .A_1       (addKernel_17_S[39:0] ), //i
    .A_2       (addKernel_18_S[39:0] ), //i
    .A_3       (addKernel_19_S[39:0] ), //i
    .A_4       (addKernel_20_S[39:0] ), //i
    .A_5       (addKernel_21_S[39:0] ), //i
    .A_6       (addKernel_22_S[39:0] ), //i
    .A_7       (addKernel_23_S[39:0] ), //i
    .A_8       (addKernel_24_S[39:0] ), //i
    .A_9       (addKernel_25_S[39:0] ), //i
    .A_10      (addKernel_26_S[39:0] ), //i
    .A_11      (addKernel_27_S[39:0] ), //i
    .A_12      (addKernel_28_S[39:0] ), //i
    .A_13      (addKernel_29_S[39:0] ), //i
    .A_14      (addKernel_30_S[39:0] ), //i
    .A_15      (addKernel_31_S[39:0] ), //i
    .S         (xAddTimes_137_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_138 (
    .A_0       (addKernel_32_S[39:0] ), //i
    .A_1       (addKernel_33_S[39:0] ), //i
    .A_2       (addKernel_34_S[39:0] ), //i
    .A_3       (addKernel_35_S[39:0] ), //i
    .A_4       (addKernel_36_S[39:0] ), //i
    .A_5       (addKernel_37_S[39:0] ), //i
    .A_6       (addKernel_38_S[39:0] ), //i
    .A_7       (addKernel_39_S[39:0] ), //i
    .A_8       (addKernel_40_S[39:0] ), //i
    .A_9       (addKernel_41_S[39:0] ), //i
    .A_10      (addKernel_42_S[39:0] ), //i
    .A_11      (addKernel_43_S[39:0] ), //i
    .A_12      (addKernel_44_S[39:0] ), //i
    .A_13      (addKernel_45_S[39:0] ), //i
    .A_14      (addKernel_46_S[39:0] ), //i
    .A_15      (addKernel_47_S[39:0] ), //i
    .S         (xAddTimes_138_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_139 (
    .A_0       (addKernel_48_S[39:0] ), //i
    .A_1       (addKernel_49_S[39:0] ), //i
    .A_2       (addKernel_50_S[39:0] ), //i
    .A_3       (addKernel_51_S[39:0] ), //i
    .A_4       (addKernel_52_S[39:0] ), //i
    .A_5       (addKernel_53_S[39:0] ), //i
    .A_6       (addKernel_54_S[39:0] ), //i
    .A_7       (addKernel_55_S[39:0] ), //i
    .A_8       (addKernel_56_S[39:0] ), //i
    .A_9       (addKernel_57_S[39:0] ), //i
    .A_10      (addKernel_58_S[39:0] ), //i
    .A_11      (addKernel_59_S[39:0] ), //i
    .A_12      (addKernel_60_S[39:0] ), //i
    .A_13      (addKernel_61_S[39:0] ), //i
    .A_14      (addKernel_62_S[39:0] ), //i
    .A_15      (addKernel_63_S[39:0] ), //i
    .S         (xAddTimes_139_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_140 (
    .A_0       (addKernel_64_S[39:0] ), //i
    .A_1       (addKernel_65_S[39:0] ), //i
    .A_2       (addKernel_66_S[39:0] ), //i
    .A_3       (addKernel_67_S[39:0] ), //i
    .A_4       (addKernel_68_S[39:0] ), //i
    .A_5       (addKernel_69_S[39:0] ), //i
    .A_6       (addKernel_70_S[39:0] ), //i
    .A_7       (addKernel_71_S[39:0] ), //i
    .A_8       (addKernel_72_S[39:0] ), //i
    .A_9       (addKernel_73_S[39:0] ), //i
    .A_10      (addKernel_74_S[39:0] ), //i
    .A_11      (addKernel_75_S[39:0] ), //i
    .A_12      (addKernel_76_S[39:0] ), //i
    .A_13      (addKernel_77_S[39:0] ), //i
    .A_14      (addKernel_78_S[39:0] ), //i
    .A_15      (addKernel_79_S[39:0] ), //i
    .S         (xAddTimes_140_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_141 (
    .A_0       (addKernel_80_S[39:0] ), //i
    .A_1       (addKernel_81_S[39:0] ), //i
    .A_2       (addKernel_82_S[39:0] ), //i
    .A_3       (addKernel_83_S[39:0] ), //i
    .A_4       (addKernel_84_S[39:0] ), //i
    .A_5       (addKernel_85_S[39:0] ), //i
    .A_6       (addKernel_86_S[39:0] ), //i
    .A_7       (addKernel_87_S[39:0] ), //i
    .A_8       (addKernel_88_S[39:0] ), //i
    .A_9       (addKernel_89_S[39:0] ), //i
    .A_10      (addKernel_90_S[39:0] ), //i
    .A_11      (addKernel_91_S[39:0] ), //i
    .A_12      (addKernel_92_S[39:0] ), //i
    .A_13      (addKernel_93_S[39:0] ), //i
    .A_14      (addKernel_94_S[39:0] ), //i
    .A_15      (addKernel_95_S[39:0] ), //i
    .S         (xAddTimes_141_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_142 (
    .A_0       (addKernel_96_S[39:0] ), //i
    .A_1       (addKernel_97_S[39:0] ), //i
    .A_2       (addKernel_98_S[39:0] ), //i
    .A_3       (addKernel_99_S[39:0] ), //i
    .A_4       (addKernel_100_S[39:0]), //i
    .A_5       (addKernel_101_S[39:0]), //i
    .A_6       (addKernel_102_S[39:0]), //i
    .A_7       (addKernel_103_S[39:0]), //i
    .A_8       (addKernel_104_S[39:0]), //i
    .A_9       (addKernel_105_S[39:0]), //i
    .A_10      (addKernel_106_S[39:0]), //i
    .A_11      (addKernel_107_S[39:0]), //i
    .A_12      (addKernel_108_S[39:0]), //i
    .A_13      (addKernel_109_S[39:0]), //i
    .A_14      (addKernel_110_S[39:0]), //i
    .A_15      (addKernel_111_S[39:0]), //i
    .S         (xAddTimes_142_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddTimes_128 xAddTimes_143 (
    .A_0       (addKernel_112_S[39:0]), //i
    .A_1       (addKernel_113_S[39:0]), //i
    .A_2       (addKernel_114_S[39:0]), //i
    .A_3       (addKernel_115_S[39:0]), //i
    .A_4       (addKernel_116_S[39:0]), //i
    .A_5       (addKernel_117_S[39:0]), //i
    .A_6       (addKernel_118_S[39:0]), //i
    .A_7       (addKernel_119_S[39:0]), //i
    .A_8       (addKernel_120_S[39:0]), //i
    .A_9       (addKernel_121_S[39:0]), //i
    .A_10      (addKernel_122_S[39:0]), //i
    .A_11      (addKernel_123_S[39:0]), //i
    .A_12      (addKernel_124_S[39:0]), //i
    .A_13      (addKernel_125_S[39:0]), //i
    .A_14      (addKernel_126_S[39:0]), //i
    .A_15      (addKernel_127_S[39:0]), //i
    .S         (xAddTimes_143_S[47:0]), //o
    .clk       (clk                  ), //i
    .reset     (reset                ), //i
    .softReset (softReset            )  //i
  );
  xAddChannelTimes xAddChannelTimes_16 (
    .A         (xAddChannelTimes_16_A[23:0]   ), //i
    .S         (xAddChannelTimes_16_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_17 (
    .A         (xAddChannelTimes_17_A[23:0]   ), //i
    .S         (xAddChannelTimes_17_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_18 (
    .A         (xAddChannelTimes_18_A[23:0]   ), //i
    .S         (xAddChannelTimes_18_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_19 (
    .A         (xAddChannelTimes_19_A[23:0]   ), //i
    .S         (xAddChannelTimes_19_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_20 (
    .A         (xAddChannelTimes_20_A[23:0]   ), //i
    .S         (xAddChannelTimes_20_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_21 (
    .A         (xAddChannelTimes_21_A[23:0]   ), //i
    .S         (xAddChannelTimes_21_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_22 (
    .A         (xAddChannelTimes_22_A[23:0]   ), //i
    .S         (xAddChannelTimes_22_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_23 (
    .A         (xAddChannelTimes_23_A[23:0]   ), //i
    .S         (xAddChannelTimes_23_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_24 (
    .A         (xAddChannelTimes_24_A[23:0]   ), //i
    .S         (xAddChannelTimes_24_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_25 (
    .A         (xAddChannelTimes_25_A[23:0]   ), //i
    .S         (xAddChannelTimes_25_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_26 (
    .A         (xAddChannelTimes_26_A[23:0]   ), //i
    .S         (xAddChannelTimes_26_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_27 (
    .A         (xAddChannelTimes_27_A[23:0]   ), //i
    .S         (xAddChannelTimes_27_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_28 (
    .A         (xAddChannelTimes_28_A[23:0]   ), //i
    .S         (xAddChannelTimes_28_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_29 (
    .A         (xAddChannelTimes_29_A[23:0]   ), //i
    .S         (xAddChannelTimes_29_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_30 (
    .A         (xAddChannelTimes_30_A[23:0]   ), //i
    .S         (xAddChannelTimes_30_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  xAddChannelTimes xAddChannelTimes_31 (
    .A         (xAddChannelTimes_31_A[23:0]   ), //i
    .S         (xAddChannelTimes_31_S[31:0]   ), //o
    .init      (convComputeCtrl_1_normPreValid), //i
    .clk       (clk                           ), //i
    .reset     (reset                         ), //i
    .softReset (softReset                     )  //i
  );
  Quan quan_1 (
    .dataIn_0     (xAddChannelTimes_16_S[31:0]       ), //i
    .dataIn_1     (xAddChannelTimes_17_S[31:0]       ), //i
    .dataIn_2     (xAddChannelTimes_18_S[31:0]       ), //i
    .dataIn_3     (xAddChannelTimes_19_S[31:0]       ), //i
    .dataIn_4     (xAddChannelTimes_20_S[31:0]       ), //i
    .dataIn_5     (xAddChannelTimes_21_S[31:0]       ), //i
    .dataIn_6     (xAddChannelTimes_22_S[31:0]       ), //i
    .dataIn_7     (xAddChannelTimes_23_S[31:0]       ), //i
    .dataIn_8     (xAddChannelTimes_24_S[31:0]       ), //i
    .dataIn_9     (xAddChannelTimes_25_S[31:0]       ), //i
    .dataIn_10    (xAddChannelTimes_26_S[31:0]       ), //i
    .dataIn_11    (xAddChannelTimes_27_S[31:0]       ), //i
    .dataIn_12    (xAddChannelTimes_28_S[31:0]       ), //i
    .dataIn_13    (xAddChannelTimes_29_S[31:0]       ), //i
    .dataIn_14    (xAddChannelTimes_30_S[31:0]       ), //i
    .dataIn_15    (xAddChannelTimes_31_S[31:0]       ), //i
    .biasIn       (loadWeight_1_biasRead_data[511:0] ), //i
    .scaleIn      (loadWeight_1_scaleRead_data[511:0]), //i
    .shiftIn      (loadWeight_1_shiftRead_data[511:0]), //i
    .zeroIn       (quanZeroData[7:0]                 ), //i
    .activationEn (enActivation                      ), //i
    .dataOut      (quan_1_dataOut[127:0]             ), //o
    .amendReg     (amendReg[31:0]                    ), //i
    .clk          (clk                               ), //i
    .reset        (reset                             ), //i
    .softReset    (softReset                         )  //i
  );
  Stride stride_1 (
    .sData_valid   (convComputeCtrl_1_mDataValid ), //i
    .sData_ready   (stride_1_sData_ready         ), //o
    .sData_payload (quan_1_dataOut[127:0]        ), //i
    .mData_valid   (stride_1_mData_valid         ), //o
    .mData_ready   (mFeatureData_ready           ), //i
    .mData_payload (stride_1_mData_payload[127:0]), //o
    .sReady        (stride_1_sReady              ), //o
    .complete      (stride_1_complete            ), //o
    .enStride      (enStride                     ), //i
    .rowNumIn      (rowNumIn[9:0]                ), //i
    .colNumIn      (colNumIn[9:0]                ), //i
    .channelOut    (channelOut[11:0]             ), //i
    .start         (startCu                      ), //i
    .last          (stride_1_last                ), //o
    .clk           (clk                          ), //i
    .reset         (reset                        ), //i
    .softReset     (softReset                    )  //i
  );
  assign sFeatureFirstLayerData_ready = channelIncr_1_sData_ready;
  always @(*) begin
    if(firstLayer) begin
      dataGenerate_1_sData_valid = channelIncr_1_mData_valid;
    end else begin
      dataGenerate_1_sData_valid = sFeatureData_valid;
    end
  end

  always @(*) begin
    if(firstLayer) begin
      channelIncr_1_mData_ready = dataGenerate_1_sData_ready;
    end else begin
      channelIncr_1_mData_ready = 1'b0;
    end
  end

  always @(*) begin
    if(firstLayer) begin
      dataGenerate_1_sData_payload = channelIncr_1_mData_payload;
    end else begin
      dataGenerate_1_sData_payload = sFeatureData_payload;
    end
  end

  always @(*) begin
    if(firstLayer) begin
      sFeatureData_ready = 1'b0;
    end else begin
      sFeatureData_ready = dataGenerate_1_sData_ready;
    end
  end

  assign sParaData_ready = loadWeight_1_sData_ready;
  assign copyWeightDone = loadWeight_1_copyWeightDone;
  assign waXpmSyncFifo_9_sCount = {1'd0, convComputeCtrl_1_sCount};
  assign waXpmSyncFifo_9_mCount = {1'd0, convComputeCtrl_1_mCount};
  assign _zz_b = _zz_b_18;
  assign _zz_b_1 = _zz_b_28;
  assign _zz_b_2 = _zz_b_38;
  assign _zz_b_3 = _zz_b_48;
  assign _zz_b_4 = _zz_b_58;
  assign _zz_b_5 = _zz_b_68;
  assign _zz_b_6 = _zz_b_78;
  assign _zz_b_7 = _zz_b_88;
  assign _zz_b_8 = _zz_b_98;
  assign dSP_1_a = loadWeight_1_weightRead_0_data[7 : 0];
  assign dSP_1_d = loadWeight_1_weightRead_0_data[135 : 128];
  assign dSP_1_b = _zz_b[7 : 0];
  assign dSP_2_a = loadWeight_1_weightRead_0_data[15 : 8];
  assign dSP_2_d = loadWeight_1_weightRead_0_data[143 : 136];
  assign dSP_2_b = _zz_b[15 : 8];
  assign dSP_3_a = loadWeight_1_weightRead_0_data[23 : 16];
  assign dSP_3_d = loadWeight_1_weightRead_0_data[151 : 144];
  assign dSP_3_b = _zz_b[23 : 16];
  assign dSP_4_a = loadWeight_1_weightRead_0_data[31 : 24];
  assign dSP_4_d = loadWeight_1_weightRead_0_data[159 : 152];
  assign dSP_4_b = _zz_b[31 : 24];
  assign dSP_5_a = loadWeight_1_weightRead_0_data[39 : 32];
  assign dSP_5_d = loadWeight_1_weightRead_0_data[167 : 160];
  assign dSP_5_b = _zz_b[39 : 32];
  assign dSP_6_a = loadWeight_1_weightRead_0_data[47 : 40];
  assign dSP_6_d = loadWeight_1_weightRead_0_data[175 : 168];
  assign dSP_6_b = _zz_b[47 : 40];
  assign dSP_7_a = loadWeight_1_weightRead_0_data[55 : 48];
  assign dSP_7_d = loadWeight_1_weightRead_0_data[183 : 176];
  assign dSP_7_b = _zz_b[55 : 48];
  assign dSP_8_a = loadWeight_1_weightRead_0_data[63 : 56];
  assign dSP_8_d = loadWeight_1_weightRead_0_data[191 : 184];
  assign dSP_8_b = _zz_b[63 : 56];
  assign dSP_9_a = loadWeight_1_weightRead_0_data[71 : 64];
  assign dSP_9_d = loadWeight_1_weightRead_0_data[199 : 192];
  assign dSP_9_b = _zz_b[71 : 64];
  assign dSP_10_a = loadWeight_1_weightRead_0_data[79 : 72];
  assign dSP_10_d = loadWeight_1_weightRead_0_data[207 : 200];
  assign dSP_10_b = _zz_b[79 : 72];
  assign dSP_11_a = loadWeight_1_weightRead_0_data[87 : 80];
  assign dSP_11_d = loadWeight_1_weightRead_0_data[215 : 208];
  assign dSP_11_b = _zz_b[87 : 80];
  assign dSP_12_a = loadWeight_1_weightRead_0_data[95 : 88];
  assign dSP_12_d = loadWeight_1_weightRead_0_data[223 : 216];
  assign dSP_12_b = _zz_b[95 : 88];
  assign dSP_13_a = loadWeight_1_weightRead_0_data[103 : 96];
  assign dSP_13_d = loadWeight_1_weightRead_0_data[231 : 224];
  assign dSP_13_b = _zz_b[103 : 96];
  assign dSP_14_a = loadWeight_1_weightRead_0_data[111 : 104];
  assign dSP_14_d = loadWeight_1_weightRead_0_data[239 : 232];
  assign dSP_14_b = _zz_b[111 : 104];
  assign dSP_15_a = loadWeight_1_weightRead_0_data[119 : 112];
  assign dSP_15_d = loadWeight_1_weightRead_0_data[247 : 240];
  assign dSP_15_b = _zz_b[119 : 112];
  assign dSP_16_a = loadWeight_1_weightRead_0_data[127 : 120];
  assign dSP_16_d = loadWeight_1_weightRead_0_data[255 : 248];
  assign dSP_16_b = _zz_b[127 : 120];
  assign dSP_17_a = loadWeight_1_weightRead_0_data[263 : 256];
  assign dSP_17_d = loadWeight_1_weightRead_0_data[391 : 384];
  assign dSP_17_b = _zz_b[7 : 0];
  assign dSP_18_a = loadWeight_1_weightRead_0_data[271 : 264];
  assign dSP_18_d = loadWeight_1_weightRead_0_data[399 : 392];
  assign dSP_18_b = _zz_b[15 : 8];
  assign dSP_19_a = loadWeight_1_weightRead_0_data[279 : 272];
  assign dSP_19_d = loadWeight_1_weightRead_0_data[407 : 400];
  assign dSP_19_b = _zz_b[23 : 16];
  assign dSP_20_a = loadWeight_1_weightRead_0_data[287 : 280];
  assign dSP_20_d = loadWeight_1_weightRead_0_data[415 : 408];
  assign dSP_20_b = _zz_b[31 : 24];
  assign dSP_21_a = loadWeight_1_weightRead_0_data[295 : 288];
  assign dSP_21_d = loadWeight_1_weightRead_0_data[423 : 416];
  assign dSP_21_b = _zz_b[39 : 32];
  assign dSP_22_a = loadWeight_1_weightRead_0_data[303 : 296];
  assign dSP_22_d = loadWeight_1_weightRead_0_data[431 : 424];
  assign dSP_22_b = _zz_b[47 : 40];
  assign dSP_23_a = loadWeight_1_weightRead_0_data[311 : 304];
  assign dSP_23_d = loadWeight_1_weightRead_0_data[439 : 432];
  assign dSP_23_b = _zz_b[55 : 48];
  assign dSP_24_a = loadWeight_1_weightRead_0_data[319 : 312];
  assign dSP_24_d = loadWeight_1_weightRead_0_data[447 : 440];
  assign dSP_24_b = _zz_b[63 : 56];
  assign dSP_25_a = loadWeight_1_weightRead_0_data[327 : 320];
  assign dSP_25_d = loadWeight_1_weightRead_0_data[455 : 448];
  assign dSP_25_b = _zz_b[71 : 64];
  assign dSP_26_a = loadWeight_1_weightRead_0_data[335 : 328];
  assign dSP_26_d = loadWeight_1_weightRead_0_data[463 : 456];
  assign dSP_26_b = _zz_b[79 : 72];
  assign dSP_27_a = loadWeight_1_weightRead_0_data[343 : 336];
  assign dSP_27_d = loadWeight_1_weightRead_0_data[471 : 464];
  assign dSP_27_b = _zz_b[87 : 80];
  assign dSP_28_a = loadWeight_1_weightRead_0_data[351 : 344];
  assign dSP_28_d = loadWeight_1_weightRead_0_data[479 : 472];
  assign dSP_28_b = _zz_b[95 : 88];
  assign dSP_29_a = loadWeight_1_weightRead_0_data[359 : 352];
  assign dSP_29_d = loadWeight_1_weightRead_0_data[487 : 480];
  assign dSP_29_b = _zz_b[103 : 96];
  assign dSP_30_a = loadWeight_1_weightRead_0_data[367 : 360];
  assign dSP_30_d = loadWeight_1_weightRead_0_data[495 : 488];
  assign dSP_30_b = _zz_b[111 : 104];
  assign dSP_31_a = loadWeight_1_weightRead_0_data[375 : 368];
  assign dSP_31_d = loadWeight_1_weightRead_0_data[503 : 496];
  assign dSP_31_b = _zz_b[119 : 112];
  assign dSP_32_a = loadWeight_1_weightRead_0_data[383 : 376];
  assign dSP_32_d = loadWeight_1_weightRead_0_data[511 : 504];
  assign dSP_32_b = _zz_b[127 : 120];
  assign dSP_33_a = loadWeight_1_weightRead_0_data[519 : 512];
  assign dSP_33_d = loadWeight_1_weightRead_0_data[647 : 640];
  assign dSP_33_b = _zz_b[7 : 0];
  assign dSP_34_a = loadWeight_1_weightRead_0_data[527 : 520];
  assign dSP_34_d = loadWeight_1_weightRead_0_data[655 : 648];
  assign dSP_34_b = _zz_b[15 : 8];
  assign dSP_35_a = loadWeight_1_weightRead_0_data[535 : 528];
  assign dSP_35_d = loadWeight_1_weightRead_0_data[663 : 656];
  assign dSP_35_b = _zz_b[23 : 16];
  assign dSP_36_a = loadWeight_1_weightRead_0_data[543 : 536];
  assign dSP_36_d = loadWeight_1_weightRead_0_data[671 : 664];
  assign dSP_36_b = _zz_b[31 : 24];
  assign dSP_37_a = loadWeight_1_weightRead_0_data[551 : 544];
  assign dSP_37_d = loadWeight_1_weightRead_0_data[679 : 672];
  assign dSP_37_b = _zz_b[39 : 32];
  assign dSP_38_a = loadWeight_1_weightRead_0_data[559 : 552];
  assign dSP_38_d = loadWeight_1_weightRead_0_data[687 : 680];
  assign dSP_38_b = _zz_b[47 : 40];
  assign dSP_39_a = loadWeight_1_weightRead_0_data[567 : 560];
  assign dSP_39_d = loadWeight_1_weightRead_0_data[695 : 688];
  assign dSP_39_b = _zz_b[55 : 48];
  assign dSP_40_a = loadWeight_1_weightRead_0_data[575 : 568];
  assign dSP_40_d = loadWeight_1_weightRead_0_data[703 : 696];
  assign dSP_40_b = _zz_b[63 : 56];
  assign dSP_41_a = loadWeight_1_weightRead_0_data[583 : 576];
  assign dSP_41_d = loadWeight_1_weightRead_0_data[711 : 704];
  assign dSP_41_b = _zz_b[71 : 64];
  assign dSP_42_a = loadWeight_1_weightRead_0_data[591 : 584];
  assign dSP_42_d = loadWeight_1_weightRead_0_data[719 : 712];
  assign dSP_42_b = _zz_b[79 : 72];
  assign dSP_43_a = loadWeight_1_weightRead_0_data[599 : 592];
  assign dSP_43_d = loadWeight_1_weightRead_0_data[727 : 720];
  assign dSP_43_b = _zz_b[87 : 80];
  assign dSP_44_a = loadWeight_1_weightRead_0_data[607 : 600];
  assign dSP_44_d = loadWeight_1_weightRead_0_data[735 : 728];
  assign dSP_44_b = _zz_b[95 : 88];
  assign dSP_45_a = loadWeight_1_weightRead_0_data[615 : 608];
  assign dSP_45_d = loadWeight_1_weightRead_0_data[743 : 736];
  assign dSP_45_b = _zz_b[103 : 96];
  assign dSP_46_a = loadWeight_1_weightRead_0_data[623 : 616];
  assign dSP_46_d = loadWeight_1_weightRead_0_data[751 : 744];
  assign dSP_46_b = _zz_b[111 : 104];
  assign dSP_47_a = loadWeight_1_weightRead_0_data[631 : 624];
  assign dSP_47_d = loadWeight_1_weightRead_0_data[759 : 752];
  assign dSP_47_b = _zz_b[119 : 112];
  assign dSP_48_a = loadWeight_1_weightRead_0_data[639 : 632];
  assign dSP_48_d = loadWeight_1_weightRead_0_data[767 : 760];
  assign dSP_48_b = _zz_b[127 : 120];
  assign dSP_49_a = loadWeight_1_weightRead_0_data[775 : 768];
  assign dSP_49_d = loadWeight_1_weightRead_0_data[903 : 896];
  assign dSP_49_b = _zz_b[7 : 0];
  assign dSP_50_a = loadWeight_1_weightRead_0_data[783 : 776];
  assign dSP_50_d = loadWeight_1_weightRead_0_data[911 : 904];
  assign dSP_50_b = _zz_b[15 : 8];
  assign dSP_51_a = loadWeight_1_weightRead_0_data[791 : 784];
  assign dSP_51_d = loadWeight_1_weightRead_0_data[919 : 912];
  assign dSP_51_b = _zz_b[23 : 16];
  assign dSP_52_a = loadWeight_1_weightRead_0_data[799 : 792];
  assign dSP_52_d = loadWeight_1_weightRead_0_data[927 : 920];
  assign dSP_52_b = _zz_b[31 : 24];
  assign dSP_53_a = loadWeight_1_weightRead_0_data[807 : 800];
  assign dSP_53_d = loadWeight_1_weightRead_0_data[935 : 928];
  assign dSP_53_b = _zz_b[39 : 32];
  assign dSP_54_a = loadWeight_1_weightRead_0_data[815 : 808];
  assign dSP_54_d = loadWeight_1_weightRead_0_data[943 : 936];
  assign dSP_54_b = _zz_b[47 : 40];
  assign dSP_55_a = loadWeight_1_weightRead_0_data[823 : 816];
  assign dSP_55_d = loadWeight_1_weightRead_0_data[951 : 944];
  assign dSP_55_b = _zz_b[55 : 48];
  assign dSP_56_a = loadWeight_1_weightRead_0_data[831 : 824];
  assign dSP_56_d = loadWeight_1_weightRead_0_data[959 : 952];
  assign dSP_56_b = _zz_b[63 : 56];
  assign dSP_57_a = loadWeight_1_weightRead_0_data[839 : 832];
  assign dSP_57_d = loadWeight_1_weightRead_0_data[967 : 960];
  assign dSP_57_b = _zz_b[71 : 64];
  assign dSP_58_a = loadWeight_1_weightRead_0_data[847 : 840];
  assign dSP_58_d = loadWeight_1_weightRead_0_data[975 : 968];
  assign dSP_58_b = _zz_b[79 : 72];
  assign dSP_59_a = loadWeight_1_weightRead_0_data[855 : 848];
  assign dSP_59_d = loadWeight_1_weightRead_0_data[983 : 976];
  assign dSP_59_b = _zz_b[87 : 80];
  assign dSP_60_a = loadWeight_1_weightRead_0_data[863 : 856];
  assign dSP_60_d = loadWeight_1_weightRead_0_data[991 : 984];
  assign dSP_60_b = _zz_b[95 : 88];
  assign dSP_61_a = loadWeight_1_weightRead_0_data[871 : 864];
  assign dSP_61_d = loadWeight_1_weightRead_0_data[999 : 992];
  assign dSP_61_b = _zz_b[103 : 96];
  assign dSP_62_a = loadWeight_1_weightRead_0_data[879 : 872];
  assign dSP_62_d = loadWeight_1_weightRead_0_data[1007 : 1000];
  assign dSP_62_b = _zz_b[111 : 104];
  assign dSP_63_a = loadWeight_1_weightRead_0_data[887 : 880];
  assign dSP_63_d = loadWeight_1_weightRead_0_data[1015 : 1008];
  assign dSP_63_b = _zz_b[119 : 112];
  assign dSP_64_a = loadWeight_1_weightRead_0_data[895 : 888];
  assign dSP_64_d = loadWeight_1_weightRead_0_data[1023 : 1016];
  assign dSP_64_b = _zz_b[127 : 120];
  assign dSP_65_a = loadWeight_1_weightRead_0_data[1031 : 1024];
  assign dSP_65_d = loadWeight_1_weightRead_0_data[1159 : 1152];
  assign dSP_65_b = _zz_b[7 : 0];
  assign dSP_66_a = loadWeight_1_weightRead_0_data[1039 : 1032];
  assign dSP_66_d = loadWeight_1_weightRead_0_data[1167 : 1160];
  assign dSP_66_b = _zz_b[15 : 8];
  assign dSP_67_a = loadWeight_1_weightRead_0_data[1047 : 1040];
  assign dSP_67_d = loadWeight_1_weightRead_0_data[1175 : 1168];
  assign dSP_67_b = _zz_b[23 : 16];
  assign dSP_68_a = loadWeight_1_weightRead_0_data[1055 : 1048];
  assign dSP_68_d = loadWeight_1_weightRead_0_data[1183 : 1176];
  assign dSP_68_b = _zz_b[31 : 24];
  assign dSP_69_a = loadWeight_1_weightRead_0_data[1063 : 1056];
  assign dSP_69_d = loadWeight_1_weightRead_0_data[1191 : 1184];
  assign dSP_69_b = _zz_b[39 : 32];
  assign dSP_70_a = loadWeight_1_weightRead_0_data[1071 : 1064];
  assign dSP_70_d = loadWeight_1_weightRead_0_data[1199 : 1192];
  assign dSP_70_b = _zz_b[47 : 40];
  assign dSP_71_a = loadWeight_1_weightRead_0_data[1079 : 1072];
  assign dSP_71_d = loadWeight_1_weightRead_0_data[1207 : 1200];
  assign dSP_71_b = _zz_b[55 : 48];
  assign dSP_72_a = loadWeight_1_weightRead_0_data[1087 : 1080];
  assign dSP_72_d = loadWeight_1_weightRead_0_data[1215 : 1208];
  assign dSP_72_b = _zz_b[63 : 56];
  assign dSP_73_a = loadWeight_1_weightRead_0_data[1095 : 1088];
  assign dSP_73_d = loadWeight_1_weightRead_0_data[1223 : 1216];
  assign dSP_73_b = _zz_b[71 : 64];
  assign dSP_74_a = loadWeight_1_weightRead_0_data[1103 : 1096];
  assign dSP_74_d = loadWeight_1_weightRead_0_data[1231 : 1224];
  assign dSP_74_b = _zz_b[79 : 72];
  assign dSP_75_a = loadWeight_1_weightRead_0_data[1111 : 1104];
  assign dSP_75_d = loadWeight_1_weightRead_0_data[1239 : 1232];
  assign dSP_75_b = _zz_b[87 : 80];
  assign dSP_76_a = loadWeight_1_weightRead_0_data[1119 : 1112];
  assign dSP_76_d = loadWeight_1_weightRead_0_data[1247 : 1240];
  assign dSP_76_b = _zz_b[95 : 88];
  assign dSP_77_a = loadWeight_1_weightRead_0_data[1127 : 1120];
  assign dSP_77_d = loadWeight_1_weightRead_0_data[1255 : 1248];
  assign dSP_77_b = _zz_b[103 : 96];
  assign dSP_78_a = loadWeight_1_weightRead_0_data[1135 : 1128];
  assign dSP_78_d = loadWeight_1_weightRead_0_data[1263 : 1256];
  assign dSP_78_b = _zz_b[111 : 104];
  assign dSP_79_a = loadWeight_1_weightRead_0_data[1143 : 1136];
  assign dSP_79_d = loadWeight_1_weightRead_0_data[1271 : 1264];
  assign dSP_79_b = _zz_b[119 : 112];
  assign dSP_80_a = loadWeight_1_weightRead_0_data[1151 : 1144];
  assign dSP_80_d = loadWeight_1_weightRead_0_data[1279 : 1272];
  assign dSP_80_b = _zz_b[127 : 120];
  assign dSP_81_a = loadWeight_1_weightRead_0_data[1287 : 1280];
  assign dSP_81_d = loadWeight_1_weightRead_0_data[1415 : 1408];
  assign dSP_81_b = _zz_b[7 : 0];
  assign dSP_82_a = loadWeight_1_weightRead_0_data[1295 : 1288];
  assign dSP_82_d = loadWeight_1_weightRead_0_data[1423 : 1416];
  assign dSP_82_b = _zz_b[15 : 8];
  assign dSP_83_a = loadWeight_1_weightRead_0_data[1303 : 1296];
  assign dSP_83_d = loadWeight_1_weightRead_0_data[1431 : 1424];
  assign dSP_83_b = _zz_b[23 : 16];
  assign dSP_84_a = loadWeight_1_weightRead_0_data[1311 : 1304];
  assign dSP_84_d = loadWeight_1_weightRead_0_data[1439 : 1432];
  assign dSP_84_b = _zz_b[31 : 24];
  assign dSP_85_a = loadWeight_1_weightRead_0_data[1319 : 1312];
  assign dSP_85_d = loadWeight_1_weightRead_0_data[1447 : 1440];
  assign dSP_85_b = _zz_b[39 : 32];
  assign dSP_86_a = loadWeight_1_weightRead_0_data[1327 : 1320];
  assign dSP_86_d = loadWeight_1_weightRead_0_data[1455 : 1448];
  assign dSP_86_b = _zz_b[47 : 40];
  assign dSP_87_a = loadWeight_1_weightRead_0_data[1335 : 1328];
  assign dSP_87_d = loadWeight_1_weightRead_0_data[1463 : 1456];
  assign dSP_87_b = _zz_b[55 : 48];
  assign dSP_88_a = loadWeight_1_weightRead_0_data[1343 : 1336];
  assign dSP_88_d = loadWeight_1_weightRead_0_data[1471 : 1464];
  assign dSP_88_b = _zz_b[63 : 56];
  assign dSP_89_a = loadWeight_1_weightRead_0_data[1351 : 1344];
  assign dSP_89_d = loadWeight_1_weightRead_0_data[1479 : 1472];
  assign dSP_89_b = _zz_b[71 : 64];
  assign dSP_90_a = loadWeight_1_weightRead_0_data[1359 : 1352];
  assign dSP_90_d = loadWeight_1_weightRead_0_data[1487 : 1480];
  assign dSP_90_b = _zz_b[79 : 72];
  assign dSP_91_a = loadWeight_1_weightRead_0_data[1367 : 1360];
  assign dSP_91_d = loadWeight_1_weightRead_0_data[1495 : 1488];
  assign dSP_91_b = _zz_b[87 : 80];
  assign dSP_92_a = loadWeight_1_weightRead_0_data[1375 : 1368];
  assign dSP_92_d = loadWeight_1_weightRead_0_data[1503 : 1496];
  assign dSP_92_b = _zz_b[95 : 88];
  assign dSP_93_a = loadWeight_1_weightRead_0_data[1383 : 1376];
  assign dSP_93_d = loadWeight_1_weightRead_0_data[1511 : 1504];
  assign dSP_93_b = _zz_b[103 : 96];
  assign dSP_94_a = loadWeight_1_weightRead_0_data[1391 : 1384];
  assign dSP_94_d = loadWeight_1_weightRead_0_data[1519 : 1512];
  assign dSP_94_b = _zz_b[111 : 104];
  assign dSP_95_a = loadWeight_1_weightRead_0_data[1399 : 1392];
  assign dSP_95_d = loadWeight_1_weightRead_0_data[1527 : 1520];
  assign dSP_95_b = _zz_b[119 : 112];
  assign dSP_96_a = loadWeight_1_weightRead_0_data[1407 : 1400];
  assign dSP_96_d = loadWeight_1_weightRead_0_data[1535 : 1528];
  assign dSP_96_b = _zz_b[127 : 120];
  assign dSP_97_a = loadWeight_1_weightRead_0_data[1543 : 1536];
  assign dSP_97_d = loadWeight_1_weightRead_0_data[1671 : 1664];
  assign dSP_97_b = _zz_b[7 : 0];
  assign dSP_98_a = loadWeight_1_weightRead_0_data[1551 : 1544];
  assign dSP_98_d = loadWeight_1_weightRead_0_data[1679 : 1672];
  assign dSP_98_b = _zz_b[15 : 8];
  assign dSP_99_a = loadWeight_1_weightRead_0_data[1559 : 1552];
  assign dSP_99_d = loadWeight_1_weightRead_0_data[1687 : 1680];
  assign dSP_99_b = _zz_b[23 : 16];
  assign dSP_100_a = loadWeight_1_weightRead_0_data[1567 : 1560];
  assign dSP_100_d = loadWeight_1_weightRead_0_data[1695 : 1688];
  assign dSP_100_b = _zz_b[31 : 24];
  assign dSP_101_a = loadWeight_1_weightRead_0_data[1575 : 1568];
  assign dSP_101_d = loadWeight_1_weightRead_0_data[1703 : 1696];
  assign dSP_101_b = _zz_b[39 : 32];
  assign dSP_102_a = loadWeight_1_weightRead_0_data[1583 : 1576];
  assign dSP_102_d = loadWeight_1_weightRead_0_data[1711 : 1704];
  assign dSP_102_b = _zz_b[47 : 40];
  assign dSP_103_a = loadWeight_1_weightRead_0_data[1591 : 1584];
  assign dSP_103_d = loadWeight_1_weightRead_0_data[1719 : 1712];
  assign dSP_103_b = _zz_b[55 : 48];
  assign dSP_104_a = loadWeight_1_weightRead_0_data[1599 : 1592];
  assign dSP_104_d = loadWeight_1_weightRead_0_data[1727 : 1720];
  assign dSP_104_b = _zz_b[63 : 56];
  assign dSP_105_a = loadWeight_1_weightRead_0_data[1607 : 1600];
  assign dSP_105_d = loadWeight_1_weightRead_0_data[1735 : 1728];
  assign dSP_105_b = _zz_b[71 : 64];
  assign dSP_106_a = loadWeight_1_weightRead_0_data[1615 : 1608];
  assign dSP_106_d = loadWeight_1_weightRead_0_data[1743 : 1736];
  assign dSP_106_b = _zz_b[79 : 72];
  assign dSP_107_a = loadWeight_1_weightRead_0_data[1623 : 1616];
  assign dSP_107_d = loadWeight_1_weightRead_0_data[1751 : 1744];
  assign dSP_107_b = _zz_b[87 : 80];
  assign dSP_108_a = loadWeight_1_weightRead_0_data[1631 : 1624];
  assign dSP_108_d = loadWeight_1_weightRead_0_data[1759 : 1752];
  assign dSP_108_b = _zz_b[95 : 88];
  assign dSP_109_a = loadWeight_1_weightRead_0_data[1639 : 1632];
  assign dSP_109_d = loadWeight_1_weightRead_0_data[1767 : 1760];
  assign dSP_109_b = _zz_b[103 : 96];
  assign dSP_110_a = loadWeight_1_weightRead_0_data[1647 : 1640];
  assign dSP_110_d = loadWeight_1_weightRead_0_data[1775 : 1768];
  assign dSP_110_b = _zz_b[111 : 104];
  assign dSP_111_a = loadWeight_1_weightRead_0_data[1655 : 1648];
  assign dSP_111_d = loadWeight_1_weightRead_0_data[1783 : 1776];
  assign dSP_111_b = _zz_b[119 : 112];
  assign dSP_112_a = loadWeight_1_weightRead_0_data[1663 : 1656];
  assign dSP_112_d = loadWeight_1_weightRead_0_data[1791 : 1784];
  assign dSP_112_b = _zz_b[127 : 120];
  assign dSP_113_a = loadWeight_1_weightRead_0_data[1799 : 1792];
  assign dSP_113_d = loadWeight_1_weightRead_0_data[1927 : 1920];
  assign dSP_113_b = _zz_b[7 : 0];
  assign dSP_114_a = loadWeight_1_weightRead_0_data[1807 : 1800];
  assign dSP_114_d = loadWeight_1_weightRead_0_data[1935 : 1928];
  assign dSP_114_b = _zz_b[15 : 8];
  assign dSP_115_a = loadWeight_1_weightRead_0_data[1815 : 1808];
  assign dSP_115_d = loadWeight_1_weightRead_0_data[1943 : 1936];
  assign dSP_115_b = _zz_b[23 : 16];
  assign dSP_116_a = loadWeight_1_weightRead_0_data[1823 : 1816];
  assign dSP_116_d = loadWeight_1_weightRead_0_data[1951 : 1944];
  assign dSP_116_b = _zz_b[31 : 24];
  assign dSP_117_a = loadWeight_1_weightRead_0_data[1831 : 1824];
  assign dSP_117_d = loadWeight_1_weightRead_0_data[1959 : 1952];
  assign dSP_117_b = _zz_b[39 : 32];
  assign dSP_118_a = loadWeight_1_weightRead_0_data[1839 : 1832];
  assign dSP_118_d = loadWeight_1_weightRead_0_data[1967 : 1960];
  assign dSP_118_b = _zz_b[47 : 40];
  assign dSP_119_a = loadWeight_1_weightRead_0_data[1847 : 1840];
  assign dSP_119_d = loadWeight_1_weightRead_0_data[1975 : 1968];
  assign dSP_119_b = _zz_b[55 : 48];
  assign dSP_120_a = loadWeight_1_weightRead_0_data[1855 : 1848];
  assign dSP_120_d = loadWeight_1_weightRead_0_data[1983 : 1976];
  assign dSP_120_b = _zz_b[63 : 56];
  assign dSP_121_a = loadWeight_1_weightRead_0_data[1863 : 1856];
  assign dSP_121_d = loadWeight_1_weightRead_0_data[1991 : 1984];
  assign dSP_121_b = _zz_b[71 : 64];
  assign dSP_122_a = loadWeight_1_weightRead_0_data[1871 : 1864];
  assign dSP_122_d = loadWeight_1_weightRead_0_data[1999 : 1992];
  assign dSP_122_b = _zz_b[79 : 72];
  assign dSP_123_a = loadWeight_1_weightRead_0_data[1879 : 1872];
  assign dSP_123_d = loadWeight_1_weightRead_0_data[2007 : 2000];
  assign dSP_123_b = _zz_b[87 : 80];
  assign dSP_124_a = loadWeight_1_weightRead_0_data[1887 : 1880];
  assign dSP_124_d = loadWeight_1_weightRead_0_data[2015 : 2008];
  assign dSP_124_b = _zz_b[95 : 88];
  assign dSP_125_a = loadWeight_1_weightRead_0_data[1895 : 1888];
  assign dSP_125_d = loadWeight_1_weightRead_0_data[2023 : 2016];
  assign dSP_125_b = _zz_b[103 : 96];
  assign dSP_126_a = loadWeight_1_weightRead_0_data[1903 : 1896];
  assign dSP_126_d = loadWeight_1_weightRead_0_data[2031 : 2024];
  assign dSP_126_b = _zz_b[111 : 104];
  assign dSP_127_a = loadWeight_1_weightRead_0_data[1911 : 1904];
  assign dSP_127_d = loadWeight_1_weightRead_0_data[2039 : 2032];
  assign dSP_127_b = _zz_b[119 : 112];
  assign dSP_128_a = loadWeight_1_weightRead_0_data[1919 : 1912];
  assign dSP_128_d = loadWeight_1_weightRead_0_data[2047 : 2040];
  assign dSP_128_b = _zz_b[127 : 120];
  assign dSP_129_a = loadWeight_1_weightRead_1_data[7 : 0];
  assign dSP_129_d = loadWeight_1_weightRead_1_data[135 : 128];
  assign dSP_129_b = _zz_b_1[7 : 0];
  assign dSP_130_a = loadWeight_1_weightRead_1_data[15 : 8];
  assign dSP_130_d = loadWeight_1_weightRead_1_data[143 : 136];
  assign dSP_130_b = _zz_b_1[15 : 8];
  assign dSP_131_a = loadWeight_1_weightRead_1_data[23 : 16];
  assign dSP_131_d = loadWeight_1_weightRead_1_data[151 : 144];
  assign dSP_131_b = _zz_b_1[23 : 16];
  assign dSP_132_a = loadWeight_1_weightRead_1_data[31 : 24];
  assign dSP_132_d = loadWeight_1_weightRead_1_data[159 : 152];
  assign dSP_132_b = _zz_b_1[31 : 24];
  assign dSP_133_a = loadWeight_1_weightRead_1_data[39 : 32];
  assign dSP_133_d = loadWeight_1_weightRead_1_data[167 : 160];
  assign dSP_133_b = _zz_b_1[39 : 32];
  assign dSP_134_a = loadWeight_1_weightRead_1_data[47 : 40];
  assign dSP_134_d = loadWeight_1_weightRead_1_data[175 : 168];
  assign dSP_134_b = _zz_b_1[47 : 40];
  assign dSP_135_a = loadWeight_1_weightRead_1_data[55 : 48];
  assign dSP_135_d = loadWeight_1_weightRead_1_data[183 : 176];
  assign dSP_135_b = _zz_b_1[55 : 48];
  assign dSP_136_a = loadWeight_1_weightRead_1_data[63 : 56];
  assign dSP_136_d = loadWeight_1_weightRead_1_data[191 : 184];
  assign dSP_136_b = _zz_b_1[63 : 56];
  assign dSP_137_a = loadWeight_1_weightRead_1_data[71 : 64];
  assign dSP_137_d = loadWeight_1_weightRead_1_data[199 : 192];
  assign dSP_137_b = _zz_b_1[71 : 64];
  assign dSP_138_a = loadWeight_1_weightRead_1_data[79 : 72];
  assign dSP_138_d = loadWeight_1_weightRead_1_data[207 : 200];
  assign dSP_138_b = _zz_b_1[79 : 72];
  assign dSP_139_a = loadWeight_1_weightRead_1_data[87 : 80];
  assign dSP_139_d = loadWeight_1_weightRead_1_data[215 : 208];
  assign dSP_139_b = _zz_b_1[87 : 80];
  assign dSP_140_a = loadWeight_1_weightRead_1_data[95 : 88];
  assign dSP_140_d = loadWeight_1_weightRead_1_data[223 : 216];
  assign dSP_140_b = _zz_b_1[95 : 88];
  assign dSP_141_a = loadWeight_1_weightRead_1_data[103 : 96];
  assign dSP_141_d = loadWeight_1_weightRead_1_data[231 : 224];
  assign dSP_141_b = _zz_b_1[103 : 96];
  assign dSP_142_a = loadWeight_1_weightRead_1_data[111 : 104];
  assign dSP_142_d = loadWeight_1_weightRead_1_data[239 : 232];
  assign dSP_142_b = _zz_b_1[111 : 104];
  assign dSP_143_a = loadWeight_1_weightRead_1_data[119 : 112];
  assign dSP_143_d = loadWeight_1_weightRead_1_data[247 : 240];
  assign dSP_143_b = _zz_b_1[119 : 112];
  assign dSP_144_a = loadWeight_1_weightRead_1_data[127 : 120];
  assign dSP_144_d = loadWeight_1_weightRead_1_data[255 : 248];
  assign dSP_144_b = _zz_b_1[127 : 120];
  assign dSP_145_a = loadWeight_1_weightRead_1_data[263 : 256];
  assign dSP_145_d = loadWeight_1_weightRead_1_data[391 : 384];
  assign dSP_145_b = _zz_b_1[7 : 0];
  assign dSP_146_a = loadWeight_1_weightRead_1_data[271 : 264];
  assign dSP_146_d = loadWeight_1_weightRead_1_data[399 : 392];
  assign dSP_146_b = _zz_b_1[15 : 8];
  assign dSP_147_a = loadWeight_1_weightRead_1_data[279 : 272];
  assign dSP_147_d = loadWeight_1_weightRead_1_data[407 : 400];
  assign dSP_147_b = _zz_b_1[23 : 16];
  assign dSP_148_a = loadWeight_1_weightRead_1_data[287 : 280];
  assign dSP_148_d = loadWeight_1_weightRead_1_data[415 : 408];
  assign dSP_148_b = _zz_b_1[31 : 24];
  assign dSP_149_a = loadWeight_1_weightRead_1_data[295 : 288];
  assign dSP_149_d = loadWeight_1_weightRead_1_data[423 : 416];
  assign dSP_149_b = _zz_b_1[39 : 32];
  assign dSP_150_a = loadWeight_1_weightRead_1_data[303 : 296];
  assign dSP_150_d = loadWeight_1_weightRead_1_data[431 : 424];
  assign dSP_150_b = _zz_b_1[47 : 40];
  assign dSP_151_a = loadWeight_1_weightRead_1_data[311 : 304];
  assign dSP_151_d = loadWeight_1_weightRead_1_data[439 : 432];
  assign dSP_151_b = _zz_b_1[55 : 48];
  assign dSP_152_a = loadWeight_1_weightRead_1_data[319 : 312];
  assign dSP_152_d = loadWeight_1_weightRead_1_data[447 : 440];
  assign dSP_152_b = _zz_b_1[63 : 56];
  assign dSP_153_a = loadWeight_1_weightRead_1_data[327 : 320];
  assign dSP_153_d = loadWeight_1_weightRead_1_data[455 : 448];
  assign dSP_153_b = _zz_b_1[71 : 64];
  assign dSP_154_a = loadWeight_1_weightRead_1_data[335 : 328];
  assign dSP_154_d = loadWeight_1_weightRead_1_data[463 : 456];
  assign dSP_154_b = _zz_b_1[79 : 72];
  assign dSP_155_a = loadWeight_1_weightRead_1_data[343 : 336];
  assign dSP_155_d = loadWeight_1_weightRead_1_data[471 : 464];
  assign dSP_155_b = _zz_b_1[87 : 80];
  assign dSP_156_a = loadWeight_1_weightRead_1_data[351 : 344];
  assign dSP_156_d = loadWeight_1_weightRead_1_data[479 : 472];
  assign dSP_156_b = _zz_b_1[95 : 88];
  assign dSP_157_a = loadWeight_1_weightRead_1_data[359 : 352];
  assign dSP_157_d = loadWeight_1_weightRead_1_data[487 : 480];
  assign dSP_157_b = _zz_b_1[103 : 96];
  assign dSP_158_a = loadWeight_1_weightRead_1_data[367 : 360];
  assign dSP_158_d = loadWeight_1_weightRead_1_data[495 : 488];
  assign dSP_158_b = _zz_b_1[111 : 104];
  assign dSP_159_a = loadWeight_1_weightRead_1_data[375 : 368];
  assign dSP_159_d = loadWeight_1_weightRead_1_data[503 : 496];
  assign dSP_159_b = _zz_b_1[119 : 112];
  assign dSP_160_a = loadWeight_1_weightRead_1_data[383 : 376];
  assign dSP_160_d = loadWeight_1_weightRead_1_data[511 : 504];
  assign dSP_160_b = _zz_b_1[127 : 120];
  assign dSP_161_a = loadWeight_1_weightRead_1_data[519 : 512];
  assign dSP_161_d = loadWeight_1_weightRead_1_data[647 : 640];
  assign dSP_161_b = _zz_b_1[7 : 0];
  assign dSP_162_a = loadWeight_1_weightRead_1_data[527 : 520];
  assign dSP_162_d = loadWeight_1_weightRead_1_data[655 : 648];
  assign dSP_162_b = _zz_b_1[15 : 8];
  assign dSP_163_a = loadWeight_1_weightRead_1_data[535 : 528];
  assign dSP_163_d = loadWeight_1_weightRead_1_data[663 : 656];
  assign dSP_163_b = _zz_b_1[23 : 16];
  assign dSP_164_a = loadWeight_1_weightRead_1_data[543 : 536];
  assign dSP_164_d = loadWeight_1_weightRead_1_data[671 : 664];
  assign dSP_164_b = _zz_b_1[31 : 24];
  assign dSP_165_a = loadWeight_1_weightRead_1_data[551 : 544];
  assign dSP_165_d = loadWeight_1_weightRead_1_data[679 : 672];
  assign dSP_165_b = _zz_b_1[39 : 32];
  assign dSP_166_a = loadWeight_1_weightRead_1_data[559 : 552];
  assign dSP_166_d = loadWeight_1_weightRead_1_data[687 : 680];
  assign dSP_166_b = _zz_b_1[47 : 40];
  assign dSP_167_a = loadWeight_1_weightRead_1_data[567 : 560];
  assign dSP_167_d = loadWeight_1_weightRead_1_data[695 : 688];
  assign dSP_167_b = _zz_b_1[55 : 48];
  assign dSP_168_a = loadWeight_1_weightRead_1_data[575 : 568];
  assign dSP_168_d = loadWeight_1_weightRead_1_data[703 : 696];
  assign dSP_168_b = _zz_b_1[63 : 56];
  assign dSP_169_a = loadWeight_1_weightRead_1_data[583 : 576];
  assign dSP_169_d = loadWeight_1_weightRead_1_data[711 : 704];
  assign dSP_169_b = _zz_b_1[71 : 64];
  assign dSP_170_a = loadWeight_1_weightRead_1_data[591 : 584];
  assign dSP_170_d = loadWeight_1_weightRead_1_data[719 : 712];
  assign dSP_170_b = _zz_b_1[79 : 72];
  assign dSP_171_a = loadWeight_1_weightRead_1_data[599 : 592];
  assign dSP_171_d = loadWeight_1_weightRead_1_data[727 : 720];
  assign dSP_171_b = _zz_b_1[87 : 80];
  assign dSP_172_a = loadWeight_1_weightRead_1_data[607 : 600];
  assign dSP_172_d = loadWeight_1_weightRead_1_data[735 : 728];
  assign dSP_172_b = _zz_b_1[95 : 88];
  assign dSP_173_a = loadWeight_1_weightRead_1_data[615 : 608];
  assign dSP_173_d = loadWeight_1_weightRead_1_data[743 : 736];
  assign dSP_173_b = _zz_b_1[103 : 96];
  assign dSP_174_a = loadWeight_1_weightRead_1_data[623 : 616];
  assign dSP_174_d = loadWeight_1_weightRead_1_data[751 : 744];
  assign dSP_174_b = _zz_b_1[111 : 104];
  assign dSP_175_a = loadWeight_1_weightRead_1_data[631 : 624];
  assign dSP_175_d = loadWeight_1_weightRead_1_data[759 : 752];
  assign dSP_175_b = _zz_b_1[119 : 112];
  assign dSP_176_a = loadWeight_1_weightRead_1_data[639 : 632];
  assign dSP_176_d = loadWeight_1_weightRead_1_data[767 : 760];
  assign dSP_176_b = _zz_b_1[127 : 120];
  assign dSP_177_a = loadWeight_1_weightRead_1_data[775 : 768];
  assign dSP_177_d = loadWeight_1_weightRead_1_data[903 : 896];
  assign dSP_177_b = _zz_b_1[7 : 0];
  assign dSP_178_a = loadWeight_1_weightRead_1_data[783 : 776];
  assign dSP_178_d = loadWeight_1_weightRead_1_data[911 : 904];
  assign dSP_178_b = _zz_b_1[15 : 8];
  assign dSP_179_a = loadWeight_1_weightRead_1_data[791 : 784];
  assign dSP_179_d = loadWeight_1_weightRead_1_data[919 : 912];
  assign dSP_179_b = _zz_b_1[23 : 16];
  assign dSP_180_a = loadWeight_1_weightRead_1_data[799 : 792];
  assign dSP_180_d = loadWeight_1_weightRead_1_data[927 : 920];
  assign dSP_180_b = _zz_b_1[31 : 24];
  assign dSP_181_a = loadWeight_1_weightRead_1_data[807 : 800];
  assign dSP_181_d = loadWeight_1_weightRead_1_data[935 : 928];
  assign dSP_181_b = _zz_b_1[39 : 32];
  assign dSP_182_a = loadWeight_1_weightRead_1_data[815 : 808];
  assign dSP_182_d = loadWeight_1_weightRead_1_data[943 : 936];
  assign dSP_182_b = _zz_b_1[47 : 40];
  assign dSP_183_a = loadWeight_1_weightRead_1_data[823 : 816];
  assign dSP_183_d = loadWeight_1_weightRead_1_data[951 : 944];
  assign dSP_183_b = _zz_b_1[55 : 48];
  assign dSP_184_a = loadWeight_1_weightRead_1_data[831 : 824];
  assign dSP_184_d = loadWeight_1_weightRead_1_data[959 : 952];
  assign dSP_184_b = _zz_b_1[63 : 56];
  assign dSP_185_a = loadWeight_1_weightRead_1_data[839 : 832];
  assign dSP_185_d = loadWeight_1_weightRead_1_data[967 : 960];
  assign dSP_185_b = _zz_b_1[71 : 64];
  assign dSP_186_a = loadWeight_1_weightRead_1_data[847 : 840];
  assign dSP_186_d = loadWeight_1_weightRead_1_data[975 : 968];
  assign dSP_186_b = _zz_b_1[79 : 72];
  assign dSP_187_a = loadWeight_1_weightRead_1_data[855 : 848];
  assign dSP_187_d = loadWeight_1_weightRead_1_data[983 : 976];
  assign dSP_187_b = _zz_b_1[87 : 80];
  assign dSP_188_a = loadWeight_1_weightRead_1_data[863 : 856];
  assign dSP_188_d = loadWeight_1_weightRead_1_data[991 : 984];
  assign dSP_188_b = _zz_b_1[95 : 88];
  assign dSP_189_a = loadWeight_1_weightRead_1_data[871 : 864];
  assign dSP_189_d = loadWeight_1_weightRead_1_data[999 : 992];
  assign dSP_189_b = _zz_b_1[103 : 96];
  assign dSP_190_a = loadWeight_1_weightRead_1_data[879 : 872];
  assign dSP_190_d = loadWeight_1_weightRead_1_data[1007 : 1000];
  assign dSP_190_b = _zz_b_1[111 : 104];
  assign dSP_191_a = loadWeight_1_weightRead_1_data[887 : 880];
  assign dSP_191_d = loadWeight_1_weightRead_1_data[1015 : 1008];
  assign dSP_191_b = _zz_b_1[119 : 112];
  assign dSP_192_a = loadWeight_1_weightRead_1_data[895 : 888];
  assign dSP_192_d = loadWeight_1_weightRead_1_data[1023 : 1016];
  assign dSP_192_b = _zz_b_1[127 : 120];
  assign dSP_193_a = loadWeight_1_weightRead_1_data[1031 : 1024];
  assign dSP_193_d = loadWeight_1_weightRead_1_data[1159 : 1152];
  assign dSP_193_b = _zz_b_1[7 : 0];
  assign dSP_194_a = loadWeight_1_weightRead_1_data[1039 : 1032];
  assign dSP_194_d = loadWeight_1_weightRead_1_data[1167 : 1160];
  assign dSP_194_b = _zz_b_1[15 : 8];
  assign dSP_195_a = loadWeight_1_weightRead_1_data[1047 : 1040];
  assign dSP_195_d = loadWeight_1_weightRead_1_data[1175 : 1168];
  assign dSP_195_b = _zz_b_1[23 : 16];
  assign dSP_196_a = loadWeight_1_weightRead_1_data[1055 : 1048];
  assign dSP_196_d = loadWeight_1_weightRead_1_data[1183 : 1176];
  assign dSP_196_b = _zz_b_1[31 : 24];
  assign dSP_197_a = loadWeight_1_weightRead_1_data[1063 : 1056];
  assign dSP_197_d = loadWeight_1_weightRead_1_data[1191 : 1184];
  assign dSP_197_b = _zz_b_1[39 : 32];
  assign dSP_198_a = loadWeight_1_weightRead_1_data[1071 : 1064];
  assign dSP_198_d = loadWeight_1_weightRead_1_data[1199 : 1192];
  assign dSP_198_b = _zz_b_1[47 : 40];
  assign dSP_199_a = loadWeight_1_weightRead_1_data[1079 : 1072];
  assign dSP_199_d = loadWeight_1_weightRead_1_data[1207 : 1200];
  assign dSP_199_b = _zz_b_1[55 : 48];
  assign dSP_200_a = loadWeight_1_weightRead_1_data[1087 : 1080];
  assign dSP_200_d = loadWeight_1_weightRead_1_data[1215 : 1208];
  assign dSP_200_b = _zz_b_1[63 : 56];
  assign dSP_201_a = loadWeight_1_weightRead_1_data[1095 : 1088];
  assign dSP_201_d = loadWeight_1_weightRead_1_data[1223 : 1216];
  assign dSP_201_b = _zz_b_1[71 : 64];
  assign dSP_202_a = loadWeight_1_weightRead_1_data[1103 : 1096];
  assign dSP_202_d = loadWeight_1_weightRead_1_data[1231 : 1224];
  assign dSP_202_b = _zz_b_1[79 : 72];
  assign dSP_203_a = loadWeight_1_weightRead_1_data[1111 : 1104];
  assign dSP_203_d = loadWeight_1_weightRead_1_data[1239 : 1232];
  assign dSP_203_b = _zz_b_1[87 : 80];
  assign dSP_204_a = loadWeight_1_weightRead_1_data[1119 : 1112];
  assign dSP_204_d = loadWeight_1_weightRead_1_data[1247 : 1240];
  assign dSP_204_b = _zz_b_1[95 : 88];
  assign dSP_205_a = loadWeight_1_weightRead_1_data[1127 : 1120];
  assign dSP_205_d = loadWeight_1_weightRead_1_data[1255 : 1248];
  assign dSP_205_b = _zz_b_1[103 : 96];
  assign dSP_206_a = loadWeight_1_weightRead_1_data[1135 : 1128];
  assign dSP_206_d = loadWeight_1_weightRead_1_data[1263 : 1256];
  assign dSP_206_b = _zz_b_1[111 : 104];
  assign dSP_207_a = loadWeight_1_weightRead_1_data[1143 : 1136];
  assign dSP_207_d = loadWeight_1_weightRead_1_data[1271 : 1264];
  assign dSP_207_b = _zz_b_1[119 : 112];
  assign dSP_208_a = loadWeight_1_weightRead_1_data[1151 : 1144];
  assign dSP_208_d = loadWeight_1_weightRead_1_data[1279 : 1272];
  assign dSP_208_b = _zz_b_1[127 : 120];
  assign dSP_209_a = loadWeight_1_weightRead_1_data[1287 : 1280];
  assign dSP_209_d = loadWeight_1_weightRead_1_data[1415 : 1408];
  assign dSP_209_b = _zz_b_1[7 : 0];
  assign dSP_210_a = loadWeight_1_weightRead_1_data[1295 : 1288];
  assign dSP_210_d = loadWeight_1_weightRead_1_data[1423 : 1416];
  assign dSP_210_b = _zz_b_1[15 : 8];
  assign dSP_211_a = loadWeight_1_weightRead_1_data[1303 : 1296];
  assign dSP_211_d = loadWeight_1_weightRead_1_data[1431 : 1424];
  assign dSP_211_b = _zz_b_1[23 : 16];
  assign dSP_212_a = loadWeight_1_weightRead_1_data[1311 : 1304];
  assign dSP_212_d = loadWeight_1_weightRead_1_data[1439 : 1432];
  assign dSP_212_b = _zz_b_1[31 : 24];
  assign dSP_213_a = loadWeight_1_weightRead_1_data[1319 : 1312];
  assign dSP_213_d = loadWeight_1_weightRead_1_data[1447 : 1440];
  assign dSP_213_b = _zz_b_1[39 : 32];
  assign dSP_214_a = loadWeight_1_weightRead_1_data[1327 : 1320];
  assign dSP_214_d = loadWeight_1_weightRead_1_data[1455 : 1448];
  assign dSP_214_b = _zz_b_1[47 : 40];
  assign dSP_215_a = loadWeight_1_weightRead_1_data[1335 : 1328];
  assign dSP_215_d = loadWeight_1_weightRead_1_data[1463 : 1456];
  assign dSP_215_b = _zz_b_1[55 : 48];
  assign dSP_216_a = loadWeight_1_weightRead_1_data[1343 : 1336];
  assign dSP_216_d = loadWeight_1_weightRead_1_data[1471 : 1464];
  assign dSP_216_b = _zz_b_1[63 : 56];
  assign dSP_217_a = loadWeight_1_weightRead_1_data[1351 : 1344];
  assign dSP_217_d = loadWeight_1_weightRead_1_data[1479 : 1472];
  assign dSP_217_b = _zz_b_1[71 : 64];
  assign dSP_218_a = loadWeight_1_weightRead_1_data[1359 : 1352];
  assign dSP_218_d = loadWeight_1_weightRead_1_data[1487 : 1480];
  assign dSP_218_b = _zz_b_1[79 : 72];
  assign dSP_219_a = loadWeight_1_weightRead_1_data[1367 : 1360];
  assign dSP_219_d = loadWeight_1_weightRead_1_data[1495 : 1488];
  assign dSP_219_b = _zz_b_1[87 : 80];
  assign dSP_220_a = loadWeight_1_weightRead_1_data[1375 : 1368];
  assign dSP_220_d = loadWeight_1_weightRead_1_data[1503 : 1496];
  assign dSP_220_b = _zz_b_1[95 : 88];
  assign dSP_221_a = loadWeight_1_weightRead_1_data[1383 : 1376];
  assign dSP_221_d = loadWeight_1_weightRead_1_data[1511 : 1504];
  assign dSP_221_b = _zz_b_1[103 : 96];
  assign dSP_222_a = loadWeight_1_weightRead_1_data[1391 : 1384];
  assign dSP_222_d = loadWeight_1_weightRead_1_data[1519 : 1512];
  assign dSP_222_b = _zz_b_1[111 : 104];
  assign dSP_223_a = loadWeight_1_weightRead_1_data[1399 : 1392];
  assign dSP_223_d = loadWeight_1_weightRead_1_data[1527 : 1520];
  assign dSP_223_b = _zz_b_1[119 : 112];
  assign dSP_224_a = loadWeight_1_weightRead_1_data[1407 : 1400];
  assign dSP_224_d = loadWeight_1_weightRead_1_data[1535 : 1528];
  assign dSP_224_b = _zz_b_1[127 : 120];
  assign dSP_225_a = loadWeight_1_weightRead_1_data[1543 : 1536];
  assign dSP_225_d = loadWeight_1_weightRead_1_data[1671 : 1664];
  assign dSP_225_b = _zz_b_1[7 : 0];
  assign dSP_226_a = loadWeight_1_weightRead_1_data[1551 : 1544];
  assign dSP_226_d = loadWeight_1_weightRead_1_data[1679 : 1672];
  assign dSP_226_b = _zz_b_1[15 : 8];
  assign dSP_227_a = loadWeight_1_weightRead_1_data[1559 : 1552];
  assign dSP_227_d = loadWeight_1_weightRead_1_data[1687 : 1680];
  assign dSP_227_b = _zz_b_1[23 : 16];
  assign dSP_228_a = loadWeight_1_weightRead_1_data[1567 : 1560];
  assign dSP_228_d = loadWeight_1_weightRead_1_data[1695 : 1688];
  assign dSP_228_b = _zz_b_1[31 : 24];
  assign dSP_229_a = loadWeight_1_weightRead_1_data[1575 : 1568];
  assign dSP_229_d = loadWeight_1_weightRead_1_data[1703 : 1696];
  assign dSP_229_b = _zz_b_1[39 : 32];
  assign dSP_230_a = loadWeight_1_weightRead_1_data[1583 : 1576];
  assign dSP_230_d = loadWeight_1_weightRead_1_data[1711 : 1704];
  assign dSP_230_b = _zz_b_1[47 : 40];
  assign dSP_231_a = loadWeight_1_weightRead_1_data[1591 : 1584];
  assign dSP_231_d = loadWeight_1_weightRead_1_data[1719 : 1712];
  assign dSP_231_b = _zz_b_1[55 : 48];
  assign dSP_232_a = loadWeight_1_weightRead_1_data[1599 : 1592];
  assign dSP_232_d = loadWeight_1_weightRead_1_data[1727 : 1720];
  assign dSP_232_b = _zz_b_1[63 : 56];
  assign dSP_233_a = loadWeight_1_weightRead_1_data[1607 : 1600];
  assign dSP_233_d = loadWeight_1_weightRead_1_data[1735 : 1728];
  assign dSP_233_b = _zz_b_1[71 : 64];
  assign dSP_234_a = loadWeight_1_weightRead_1_data[1615 : 1608];
  assign dSP_234_d = loadWeight_1_weightRead_1_data[1743 : 1736];
  assign dSP_234_b = _zz_b_1[79 : 72];
  assign dSP_235_a = loadWeight_1_weightRead_1_data[1623 : 1616];
  assign dSP_235_d = loadWeight_1_weightRead_1_data[1751 : 1744];
  assign dSP_235_b = _zz_b_1[87 : 80];
  assign dSP_236_a = loadWeight_1_weightRead_1_data[1631 : 1624];
  assign dSP_236_d = loadWeight_1_weightRead_1_data[1759 : 1752];
  assign dSP_236_b = _zz_b_1[95 : 88];
  assign dSP_237_a = loadWeight_1_weightRead_1_data[1639 : 1632];
  assign dSP_237_d = loadWeight_1_weightRead_1_data[1767 : 1760];
  assign dSP_237_b = _zz_b_1[103 : 96];
  assign dSP_238_a = loadWeight_1_weightRead_1_data[1647 : 1640];
  assign dSP_238_d = loadWeight_1_weightRead_1_data[1775 : 1768];
  assign dSP_238_b = _zz_b_1[111 : 104];
  assign dSP_239_a = loadWeight_1_weightRead_1_data[1655 : 1648];
  assign dSP_239_d = loadWeight_1_weightRead_1_data[1783 : 1776];
  assign dSP_239_b = _zz_b_1[119 : 112];
  assign dSP_240_a = loadWeight_1_weightRead_1_data[1663 : 1656];
  assign dSP_240_d = loadWeight_1_weightRead_1_data[1791 : 1784];
  assign dSP_240_b = _zz_b_1[127 : 120];
  assign dSP_241_a = loadWeight_1_weightRead_1_data[1799 : 1792];
  assign dSP_241_d = loadWeight_1_weightRead_1_data[1927 : 1920];
  assign dSP_241_b = _zz_b_1[7 : 0];
  assign dSP_242_a = loadWeight_1_weightRead_1_data[1807 : 1800];
  assign dSP_242_d = loadWeight_1_weightRead_1_data[1935 : 1928];
  assign dSP_242_b = _zz_b_1[15 : 8];
  assign dSP_243_a = loadWeight_1_weightRead_1_data[1815 : 1808];
  assign dSP_243_d = loadWeight_1_weightRead_1_data[1943 : 1936];
  assign dSP_243_b = _zz_b_1[23 : 16];
  assign dSP_244_a = loadWeight_1_weightRead_1_data[1823 : 1816];
  assign dSP_244_d = loadWeight_1_weightRead_1_data[1951 : 1944];
  assign dSP_244_b = _zz_b_1[31 : 24];
  assign dSP_245_a = loadWeight_1_weightRead_1_data[1831 : 1824];
  assign dSP_245_d = loadWeight_1_weightRead_1_data[1959 : 1952];
  assign dSP_245_b = _zz_b_1[39 : 32];
  assign dSP_246_a = loadWeight_1_weightRead_1_data[1839 : 1832];
  assign dSP_246_d = loadWeight_1_weightRead_1_data[1967 : 1960];
  assign dSP_246_b = _zz_b_1[47 : 40];
  assign dSP_247_a = loadWeight_1_weightRead_1_data[1847 : 1840];
  assign dSP_247_d = loadWeight_1_weightRead_1_data[1975 : 1968];
  assign dSP_247_b = _zz_b_1[55 : 48];
  assign dSP_248_a = loadWeight_1_weightRead_1_data[1855 : 1848];
  assign dSP_248_d = loadWeight_1_weightRead_1_data[1983 : 1976];
  assign dSP_248_b = _zz_b_1[63 : 56];
  assign dSP_249_a = loadWeight_1_weightRead_1_data[1863 : 1856];
  assign dSP_249_d = loadWeight_1_weightRead_1_data[1991 : 1984];
  assign dSP_249_b = _zz_b_1[71 : 64];
  assign dSP_250_a = loadWeight_1_weightRead_1_data[1871 : 1864];
  assign dSP_250_d = loadWeight_1_weightRead_1_data[1999 : 1992];
  assign dSP_250_b = _zz_b_1[79 : 72];
  assign dSP_251_a = loadWeight_1_weightRead_1_data[1879 : 1872];
  assign dSP_251_d = loadWeight_1_weightRead_1_data[2007 : 2000];
  assign dSP_251_b = _zz_b_1[87 : 80];
  assign dSP_252_a = loadWeight_1_weightRead_1_data[1887 : 1880];
  assign dSP_252_d = loadWeight_1_weightRead_1_data[2015 : 2008];
  assign dSP_252_b = _zz_b_1[95 : 88];
  assign dSP_253_a = loadWeight_1_weightRead_1_data[1895 : 1888];
  assign dSP_253_d = loadWeight_1_weightRead_1_data[2023 : 2016];
  assign dSP_253_b = _zz_b_1[103 : 96];
  assign dSP_254_a = loadWeight_1_weightRead_1_data[1903 : 1896];
  assign dSP_254_d = loadWeight_1_weightRead_1_data[2031 : 2024];
  assign dSP_254_b = _zz_b_1[111 : 104];
  assign dSP_255_a = loadWeight_1_weightRead_1_data[1911 : 1904];
  assign dSP_255_d = loadWeight_1_weightRead_1_data[2039 : 2032];
  assign dSP_255_b = _zz_b_1[119 : 112];
  assign dSP_256_a = loadWeight_1_weightRead_1_data[1919 : 1912];
  assign dSP_256_d = loadWeight_1_weightRead_1_data[2047 : 2040];
  assign dSP_256_b = _zz_b_1[127 : 120];
  assign dSP_257_a = loadWeight_1_weightRead_2_data[7 : 0];
  assign dSP_257_d = loadWeight_1_weightRead_2_data[135 : 128];
  assign dSP_257_b = _zz_b_2[7 : 0];
  assign dSP_258_a = loadWeight_1_weightRead_2_data[15 : 8];
  assign dSP_258_d = loadWeight_1_weightRead_2_data[143 : 136];
  assign dSP_258_b = _zz_b_2[15 : 8];
  assign dSP_259_a = loadWeight_1_weightRead_2_data[23 : 16];
  assign dSP_259_d = loadWeight_1_weightRead_2_data[151 : 144];
  assign dSP_259_b = _zz_b_2[23 : 16];
  assign dSP_260_a = loadWeight_1_weightRead_2_data[31 : 24];
  assign dSP_260_d = loadWeight_1_weightRead_2_data[159 : 152];
  assign dSP_260_b = _zz_b_2[31 : 24];
  assign dSP_261_a = loadWeight_1_weightRead_2_data[39 : 32];
  assign dSP_261_d = loadWeight_1_weightRead_2_data[167 : 160];
  assign dSP_261_b = _zz_b_2[39 : 32];
  assign dSP_262_a = loadWeight_1_weightRead_2_data[47 : 40];
  assign dSP_262_d = loadWeight_1_weightRead_2_data[175 : 168];
  assign dSP_262_b = _zz_b_2[47 : 40];
  assign dSP_263_a = loadWeight_1_weightRead_2_data[55 : 48];
  assign dSP_263_d = loadWeight_1_weightRead_2_data[183 : 176];
  assign dSP_263_b = _zz_b_2[55 : 48];
  assign dSP_264_a = loadWeight_1_weightRead_2_data[63 : 56];
  assign dSP_264_d = loadWeight_1_weightRead_2_data[191 : 184];
  assign dSP_264_b = _zz_b_2[63 : 56];
  assign dSP_265_a = loadWeight_1_weightRead_2_data[71 : 64];
  assign dSP_265_d = loadWeight_1_weightRead_2_data[199 : 192];
  assign dSP_265_b = _zz_b_2[71 : 64];
  assign dSP_266_a = loadWeight_1_weightRead_2_data[79 : 72];
  assign dSP_266_d = loadWeight_1_weightRead_2_data[207 : 200];
  assign dSP_266_b = _zz_b_2[79 : 72];
  assign dSP_267_a = loadWeight_1_weightRead_2_data[87 : 80];
  assign dSP_267_d = loadWeight_1_weightRead_2_data[215 : 208];
  assign dSP_267_b = _zz_b_2[87 : 80];
  assign dSP_268_a = loadWeight_1_weightRead_2_data[95 : 88];
  assign dSP_268_d = loadWeight_1_weightRead_2_data[223 : 216];
  assign dSP_268_b = _zz_b_2[95 : 88];
  assign dSP_269_a = loadWeight_1_weightRead_2_data[103 : 96];
  assign dSP_269_d = loadWeight_1_weightRead_2_data[231 : 224];
  assign dSP_269_b = _zz_b_2[103 : 96];
  assign dSP_270_a = loadWeight_1_weightRead_2_data[111 : 104];
  assign dSP_270_d = loadWeight_1_weightRead_2_data[239 : 232];
  assign dSP_270_b = _zz_b_2[111 : 104];
  assign dSP_271_a = loadWeight_1_weightRead_2_data[119 : 112];
  assign dSP_271_d = loadWeight_1_weightRead_2_data[247 : 240];
  assign dSP_271_b = _zz_b_2[119 : 112];
  assign dSP_272_a = loadWeight_1_weightRead_2_data[127 : 120];
  assign dSP_272_d = loadWeight_1_weightRead_2_data[255 : 248];
  assign dSP_272_b = _zz_b_2[127 : 120];
  assign dSP_273_a = loadWeight_1_weightRead_2_data[263 : 256];
  assign dSP_273_d = loadWeight_1_weightRead_2_data[391 : 384];
  assign dSP_273_b = _zz_b_2[7 : 0];
  assign dSP_274_a = loadWeight_1_weightRead_2_data[271 : 264];
  assign dSP_274_d = loadWeight_1_weightRead_2_data[399 : 392];
  assign dSP_274_b = _zz_b_2[15 : 8];
  assign dSP_275_a = loadWeight_1_weightRead_2_data[279 : 272];
  assign dSP_275_d = loadWeight_1_weightRead_2_data[407 : 400];
  assign dSP_275_b = _zz_b_2[23 : 16];
  assign dSP_276_a = loadWeight_1_weightRead_2_data[287 : 280];
  assign dSP_276_d = loadWeight_1_weightRead_2_data[415 : 408];
  assign dSP_276_b = _zz_b_2[31 : 24];
  assign dSP_277_a = loadWeight_1_weightRead_2_data[295 : 288];
  assign dSP_277_d = loadWeight_1_weightRead_2_data[423 : 416];
  assign dSP_277_b = _zz_b_2[39 : 32];
  assign dSP_278_a = loadWeight_1_weightRead_2_data[303 : 296];
  assign dSP_278_d = loadWeight_1_weightRead_2_data[431 : 424];
  assign dSP_278_b = _zz_b_2[47 : 40];
  assign dSP_279_a = loadWeight_1_weightRead_2_data[311 : 304];
  assign dSP_279_d = loadWeight_1_weightRead_2_data[439 : 432];
  assign dSP_279_b = _zz_b_2[55 : 48];
  assign dSP_280_a = loadWeight_1_weightRead_2_data[319 : 312];
  assign dSP_280_d = loadWeight_1_weightRead_2_data[447 : 440];
  assign dSP_280_b = _zz_b_2[63 : 56];
  assign dSP_281_a = loadWeight_1_weightRead_2_data[327 : 320];
  assign dSP_281_d = loadWeight_1_weightRead_2_data[455 : 448];
  assign dSP_281_b = _zz_b_2[71 : 64];
  assign dSP_282_a = loadWeight_1_weightRead_2_data[335 : 328];
  assign dSP_282_d = loadWeight_1_weightRead_2_data[463 : 456];
  assign dSP_282_b = _zz_b_2[79 : 72];
  assign dSP_283_a = loadWeight_1_weightRead_2_data[343 : 336];
  assign dSP_283_d = loadWeight_1_weightRead_2_data[471 : 464];
  assign dSP_283_b = _zz_b_2[87 : 80];
  assign dSP_284_a = loadWeight_1_weightRead_2_data[351 : 344];
  assign dSP_284_d = loadWeight_1_weightRead_2_data[479 : 472];
  assign dSP_284_b = _zz_b_2[95 : 88];
  assign dSP_285_a = loadWeight_1_weightRead_2_data[359 : 352];
  assign dSP_285_d = loadWeight_1_weightRead_2_data[487 : 480];
  assign dSP_285_b = _zz_b_2[103 : 96];
  assign dSP_286_a = loadWeight_1_weightRead_2_data[367 : 360];
  assign dSP_286_d = loadWeight_1_weightRead_2_data[495 : 488];
  assign dSP_286_b = _zz_b_2[111 : 104];
  assign dSP_287_a = loadWeight_1_weightRead_2_data[375 : 368];
  assign dSP_287_d = loadWeight_1_weightRead_2_data[503 : 496];
  assign dSP_287_b = _zz_b_2[119 : 112];
  assign dSP_288_a = loadWeight_1_weightRead_2_data[383 : 376];
  assign dSP_288_d = loadWeight_1_weightRead_2_data[511 : 504];
  assign dSP_288_b = _zz_b_2[127 : 120];
  assign dSP_289_a = loadWeight_1_weightRead_2_data[519 : 512];
  assign dSP_289_d = loadWeight_1_weightRead_2_data[647 : 640];
  assign dSP_289_b = _zz_b_2[7 : 0];
  assign dSP_290_a = loadWeight_1_weightRead_2_data[527 : 520];
  assign dSP_290_d = loadWeight_1_weightRead_2_data[655 : 648];
  assign dSP_290_b = _zz_b_2[15 : 8];
  assign dSP_291_a = loadWeight_1_weightRead_2_data[535 : 528];
  assign dSP_291_d = loadWeight_1_weightRead_2_data[663 : 656];
  assign dSP_291_b = _zz_b_2[23 : 16];
  assign dSP_292_a = loadWeight_1_weightRead_2_data[543 : 536];
  assign dSP_292_d = loadWeight_1_weightRead_2_data[671 : 664];
  assign dSP_292_b = _zz_b_2[31 : 24];
  assign dSP_293_a = loadWeight_1_weightRead_2_data[551 : 544];
  assign dSP_293_d = loadWeight_1_weightRead_2_data[679 : 672];
  assign dSP_293_b = _zz_b_2[39 : 32];
  assign dSP_294_a = loadWeight_1_weightRead_2_data[559 : 552];
  assign dSP_294_d = loadWeight_1_weightRead_2_data[687 : 680];
  assign dSP_294_b = _zz_b_2[47 : 40];
  assign dSP_295_a = loadWeight_1_weightRead_2_data[567 : 560];
  assign dSP_295_d = loadWeight_1_weightRead_2_data[695 : 688];
  assign dSP_295_b = _zz_b_2[55 : 48];
  assign dSP_296_a = loadWeight_1_weightRead_2_data[575 : 568];
  assign dSP_296_d = loadWeight_1_weightRead_2_data[703 : 696];
  assign dSP_296_b = _zz_b_2[63 : 56];
  assign dSP_297_a = loadWeight_1_weightRead_2_data[583 : 576];
  assign dSP_297_d = loadWeight_1_weightRead_2_data[711 : 704];
  assign dSP_297_b = _zz_b_2[71 : 64];
  assign dSP_298_a = loadWeight_1_weightRead_2_data[591 : 584];
  assign dSP_298_d = loadWeight_1_weightRead_2_data[719 : 712];
  assign dSP_298_b = _zz_b_2[79 : 72];
  assign dSP_299_a = loadWeight_1_weightRead_2_data[599 : 592];
  assign dSP_299_d = loadWeight_1_weightRead_2_data[727 : 720];
  assign dSP_299_b = _zz_b_2[87 : 80];
  assign dSP_300_a = loadWeight_1_weightRead_2_data[607 : 600];
  assign dSP_300_d = loadWeight_1_weightRead_2_data[735 : 728];
  assign dSP_300_b = _zz_b_2[95 : 88];
  assign dSP_301_a = loadWeight_1_weightRead_2_data[615 : 608];
  assign dSP_301_d = loadWeight_1_weightRead_2_data[743 : 736];
  assign dSP_301_b = _zz_b_2[103 : 96];
  assign dSP_302_a = loadWeight_1_weightRead_2_data[623 : 616];
  assign dSP_302_d = loadWeight_1_weightRead_2_data[751 : 744];
  assign dSP_302_b = _zz_b_2[111 : 104];
  assign dSP_303_a = loadWeight_1_weightRead_2_data[631 : 624];
  assign dSP_303_d = loadWeight_1_weightRead_2_data[759 : 752];
  assign dSP_303_b = _zz_b_2[119 : 112];
  assign dSP_304_a = loadWeight_1_weightRead_2_data[639 : 632];
  assign dSP_304_d = loadWeight_1_weightRead_2_data[767 : 760];
  assign dSP_304_b = _zz_b_2[127 : 120];
  assign dSP_305_a = loadWeight_1_weightRead_2_data[775 : 768];
  assign dSP_305_d = loadWeight_1_weightRead_2_data[903 : 896];
  assign dSP_305_b = _zz_b_2[7 : 0];
  assign dSP_306_a = loadWeight_1_weightRead_2_data[783 : 776];
  assign dSP_306_d = loadWeight_1_weightRead_2_data[911 : 904];
  assign dSP_306_b = _zz_b_2[15 : 8];
  assign dSP_307_a = loadWeight_1_weightRead_2_data[791 : 784];
  assign dSP_307_d = loadWeight_1_weightRead_2_data[919 : 912];
  assign dSP_307_b = _zz_b_2[23 : 16];
  assign dSP_308_a = loadWeight_1_weightRead_2_data[799 : 792];
  assign dSP_308_d = loadWeight_1_weightRead_2_data[927 : 920];
  assign dSP_308_b = _zz_b_2[31 : 24];
  assign dSP_309_a = loadWeight_1_weightRead_2_data[807 : 800];
  assign dSP_309_d = loadWeight_1_weightRead_2_data[935 : 928];
  assign dSP_309_b = _zz_b_2[39 : 32];
  assign dSP_310_a = loadWeight_1_weightRead_2_data[815 : 808];
  assign dSP_310_d = loadWeight_1_weightRead_2_data[943 : 936];
  assign dSP_310_b = _zz_b_2[47 : 40];
  assign dSP_311_a = loadWeight_1_weightRead_2_data[823 : 816];
  assign dSP_311_d = loadWeight_1_weightRead_2_data[951 : 944];
  assign dSP_311_b = _zz_b_2[55 : 48];
  assign dSP_312_a = loadWeight_1_weightRead_2_data[831 : 824];
  assign dSP_312_d = loadWeight_1_weightRead_2_data[959 : 952];
  assign dSP_312_b = _zz_b_2[63 : 56];
  assign dSP_313_a = loadWeight_1_weightRead_2_data[839 : 832];
  assign dSP_313_d = loadWeight_1_weightRead_2_data[967 : 960];
  assign dSP_313_b = _zz_b_2[71 : 64];
  assign dSP_314_a = loadWeight_1_weightRead_2_data[847 : 840];
  assign dSP_314_d = loadWeight_1_weightRead_2_data[975 : 968];
  assign dSP_314_b = _zz_b_2[79 : 72];
  assign dSP_315_a = loadWeight_1_weightRead_2_data[855 : 848];
  assign dSP_315_d = loadWeight_1_weightRead_2_data[983 : 976];
  assign dSP_315_b = _zz_b_2[87 : 80];
  assign dSP_316_a = loadWeight_1_weightRead_2_data[863 : 856];
  assign dSP_316_d = loadWeight_1_weightRead_2_data[991 : 984];
  assign dSP_316_b = _zz_b_2[95 : 88];
  assign dSP_317_a = loadWeight_1_weightRead_2_data[871 : 864];
  assign dSP_317_d = loadWeight_1_weightRead_2_data[999 : 992];
  assign dSP_317_b = _zz_b_2[103 : 96];
  assign dSP_318_a = loadWeight_1_weightRead_2_data[879 : 872];
  assign dSP_318_d = loadWeight_1_weightRead_2_data[1007 : 1000];
  assign dSP_318_b = _zz_b_2[111 : 104];
  assign dSP_319_a = loadWeight_1_weightRead_2_data[887 : 880];
  assign dSP_319_d = loadWeight_1_weightRead_2_data[1015 : 1008];
  assign dSP_319_b = _zz_b_2[119 : 112];
  assign dSP_320_a = loadWeight_1_weightRead_2_data[895 : 888];
  assign dSP_320_d = loadWeight_1_weightRead_2_data[1023 : 1016];
  assign dSP_320_b = _zz_b_2[127 : 120];
  assign dSP_321_a = loadWeight_1_weightRead_2_data[1031 : 1024];
  assign dSP_321_d = loadWeight_1_weightRead_2_data[1159 : 1152];
  assign dSP_321_b = _zz_b_2[7 : 0];
  assign dSP_322_a = loadWeight_1_weightRead_2_data[1039 : 1032];
  assign dSP_322_d = loadWeight_1_weightRead_2_data[1167 : 1160];
  assign dSP_322_b = _zz_b_2[15 : 8];
  assign dSP_323_a = loadWeight_1_weightRead_2_data[1047 : 1040];
  assign dSP_323_d = loadWeight_1_weightRead_2_data[1175 : 1168];
  assign dSP_323_b = _zz_b_2[23 : 16];
  assign dSP_324_a = loadWeight_1_weightRead_2_data[1055 : 1048];
  assign dSP_324_d = loadWeight_1_weightRead_2_data[1183 : 1176];
  assign dSP_324_b = _zz_b_2[31 : 24];
  assign dSP_325_a = loadWeight_1_weightRead_2_data[1063 : 1056];
  assign dSP_325_d = loadWeight_1_weightRead_2_data[1191 : 1184];
  assign dSP_325_b = _zz_b_2[39 : 32];
  assign dSP_326_a = loadWeight_1_weightRead_2_data[1071 : 1064];
  assign dSP_326_d = loadWeight_1_weightRead_2_data[1199 : 1192];
  assign dSP_326_b = _zz_b_2[47 : 40];
  assign dSP_327_a = loadWeight_1_weightRead_2_data[1079 : 1072];
  assign dSP_327_d = loadWeight_1_weightRead_2_data[1207 : 1200];
  assign dSP_327_b = _zz_b_2[55 : 48];
  assign dSP_328_a = loadWeight_1_weightRead_2_data[1087 : 1080];
  assign dSP_328_d = loadWeight_1_weightRead_2_data[1215 : 1208];
  assign dSP_328_b = _zz_b_2[63 : 56];
  assign dSP_329_a = loadWeight_1_weightRead_2_data[1095 : 1088];
  assign dSP_329_d = loadWeight_1_weightRead_2_data[1223 : 1216];
  assign dSP_329_b = _zz_b_2[71 : 64];
  assign dSP_330_a = loadWeight_1_weightRead_2_data[1103 : 1096];
  assign dSP_330_d = loadWeight_1_weightRead_2_data[1231 : 1224];
  assign dSP_330_b = _zz_b_2[79 : 72];
  assign dSP_331_a = loadWeight_1_weightRead_2_data[1111 : 1104];
  assign dSP_331_d = loadWeight_1_weightRead_2_data[1239 : 1232];
  assign dSP_331_b = _zz_b_2[87 : 80];
  assign dSP_332_a = loadWeight_1_weightRead_2_data[1119 : 1112];
  assign dSP_332_d = loadWeight_1_weightRead_2_data[1247 : 1240];
  assign dSP_332_b = _zz_b_2[95 : 88];
  assign dSP_333_a = loadWeight_1_weightRead_2_data[1127 : 1120];
  assign dSP_333_d = loadWeight_1_weightRead_2_data[1255 : 1248];
  assign dSP_333_b = _zz_b_2[103 : 96];
  assign dSP_334_a = loadWeight_1_weightRead_2_data[1135 : 1128];
  assign dSP_334_d = loadWeight_1_weightRead_2_data[1263 : 1256];
  assign dSP_334_b = _zz_b_2[111 : 104];
  assign dSP_335_a = loadWeight_1_weightRead_2_data[1143 : 1136];
  assign dSP_335_d = loadWeight_1_weightRead_2_data[1271 : 1264];
  assign dSP_335_b = _zz_b_2[119 : 112];
  assign dSP_336_a = loadWeight_1_weightRead_2_data[1151 : 1144];
  assign dSP_336_d = loadWeight_1_weightRead_2_data[1279 : 1272];
  assign dSP_336_b = _zz_b_2[127 : 120];
  assign dSP_337_a = loadWeight_1_weightRead_2_data[1287 : 1280];
  assign dSP_337_d = loadWeight_1_weightRead_2_data[1415 : 1408];
  assign dSP_337_b = _zz_b_2[7 : 0];
  assign dSP_338_a = loadWeight_1_weightRead_2_data[1295 : 1288];
  assign dSP_338_d = loadWeight_1_weightRead_2_data[1423 : 1416];
  assign dSP_338_b = _zz_b_2[15 : 8];
  assign dSP_339_a = loadWeight_1_weightRead_2_data[1303 : 1296];
  assign dSP_339_d = loadWeight_1_weightRead_2_data[1431 : 1424];
  assign dSP_339_b = _zz_b_2[23 : 16];
  assign dSP_340_a = loadWeight_1_weightRead_2_data[1311 : 1304];
  assign dSP_340_d = loadWeight_1_weightRead_2_data[1439 : 1432];
  assign dSP_340_b = _zz_b_2[31 : 24];
  assign dSP_341_a = loadWeight_1_weightRead_2_data[1319 : 1312];
  assign dSP_341_d = loadWeight_1_weightRead_2_data[1447 : 1440];
  assign dSP_341_b = _zz_b_2[39 : 32];
  assign dSP_342_a = loadWeight_1_weightRead_2_data[1327 : 1320];
  assign dSP_342_d = loadWeight_1_weightRead_2_data[1455 : 1448];
  assign dSP_342_b = _zz_b_2[47 : 40];
  assign dSP_343_a = loadWeight_1_weightRead_2_data[1335 : 1328];
  assign dSP_343_d = loadWeight_1_weightRead_2_data[1463 : 1456];
  assign dSP_343_b = _zz_b_2[55 : 48];
  assign dSP_344_a = loadWeight_1_weightRead_2_data[1343 : 1336];
  assign dSP_344_d = loadWeight_1_weightRead_2_data[1471 : 1464];
  assign dSP_344_b = _zz_b_2[63 : 56];
  assign dSP_345_a = loadWeight_1_weightRead_2_data[1351 : 1344];
  assign dSP_345_d = loadWeight_1_weightRead_2_data[1479 : 1472];
  assign dSP_345_b = _zz_b_2[71 : 64];
  assign dSP_346_a = loadWeight_1_weightRead_2_data[1359 : 1352];
  assign dSP_346_d = loadWeight_1_weightRead_2_data[1487 : 1480];
  assign dSP_346_b = _zz_b_2[79 : 72];
  assign dSP_347_a = loadWeight_1_weightRead_2_data[1367 : 1360];
  assign dSP_347_d = loadWeight_1_weightRead_2_data[1495 : 1488];
  assign dSP_347_b = _zz_b_2[87 : 80];
  assign dSP_348_a = loadWeight_1_weightRead_2_data[1375 : 1368];
  assign dSP_348_d = loadWeight_1_weightRead_2_data[1503 : 1496];
  assign dSP_348_b = _zz_b_2[95 : 88];
  assign dSP_349_a = loadWeight_1_weightRead_2_data[1383 : 1376];
  assign dSP_349_d = loadWeight_1_weightRead_2_data[1511 : 1504];
  assign dSP_349_b = _zz_b_2[103 : 96];
  assign dSP_350_a = loadWeight_1_weightRead_2_data[1391 : 1384];
  assign dSP_350_d = loadWeight_1_weightRead_2_data[1519 : 1512];
  assign dSP_350_b = _zz_b_2[111 : 104];
  assign dSP_351_a = loadWeight_1_weightRead_2_data[1399 : 1392];
  assign dSP_351_d = loadWeight_1_weightRead_2_data[1527 : 1520];
  assign dSP_351_b = _zz_b_2[119 : 112];
  assign dSP_352_a = loadWeight_1_weightRead_2_data[1407 : 1400];
  assign dSP_352_d = loadWeight_1_weightRead_2_data[1535 : 1528];
  assign dSP_352_b = _zz_b_2[127 : 120];
  assign dSP_353_a = loadWeight_1_weightRead_2_data[1543 : 1536];
  assign dSP_353_d = loadWeight_1_weightRead_2_data[1671 : 1664];
  assign dSP_353_b = _zz_b_2[7 : 0];
  assign dSP_354_a = loadWeight_1_weightRead_2_data[1551 : 1544];
  assign dSP_354_d = loadWeight_1_weightRead_2_data[1679 : 1672];
  assign dSP_354_b = _zz_b_2[15 : 8];
  assign dSP_355_a = loadWeight_1_weightRead_2_data[1559 : 1552];
  assign dSP_355_d = loadWeight_1_weightRead_2_data[1687 : 1680];
  assign dSP_355_b = _zz_b_2[23 : 16];
  assign dSP_356_a = loadWeight_1_weightRead_2_data[1567 : 1560];
  assign dSP_356_d = loadWeight_1_weightRead_2_data[1695 : 1688];
  assign dSP_356_b = _zz_b_2[31 : 24];
  assign dSP_357_a = loadWeight_1_weightRead_2_data[1575 : 1568];
  assign dSP_357_d = loadWeight_1_weightRead_2_data[1703 : 1696];
  assign dSP_357_b = _zz_b_2[39 : 32];
  assign dSP_358_a = loadWeight_1_weightRead_2_data[1583 : 1576];
  assign dSP_358_d = loadWeight_1_weightRead_2_data[1711 : 1704];
  assign dSP_358_b = _zz_b_2[47 : 40];
  assign dSP_359_a = loadWeight_1_weightRead_2_data[1591 : 1584];
  assign dSP_359_d = loadWeight_1_weightRead_2_data[1719 : 1712];
  assign dSP_359_b = _zz_b_2[55 : 48];
  assign dSP_360_a = loadWeight_1_weightRead_2_data[1599 : 1592];
  assign dSP_360_d = loadWeight_1_weightRead_2_data[1727 : 1720];
  assign dSP_360_b = _zz_b_2[63 : 56];
  assign dSP_361_a = loadWeight_1_weightRead_2_data[1607 : 1600];
  assign dSP_361_d = loadWeight_1_weightRead_2_data[1735 : 1728];
  assign dSP_361_b = _zz_b_2[71 : 64];
  assign dSP_362_a = loadWeight_1_weightRead_2_data[1615 : 1608];
  assign dSP_362_d = loadWeight_1_weightRead_2_data[1743 : 1736];
  assign dSP_362_b = _zz_b_2[79 : 72];
  assign dSP_363_a = loadWeight_1_weightRead_2_data[1623 : 1616];
  assign dSP_363_d = loadWeight_1_weightRead_2_data[1751 : 1744];
  assign dSP_363_b = _zz_b_2[87 : 80];
  assign dSP_364_a = loadWeight_1_weightRead_2_data[1631 : 1624];
  assign dSP_364_d = loadWeight_1_weightRead_2_data[1759 : 1752];
  assign dSP_364_b = _zz_b_2[95 : 88];
  assign dSP_365_a = loadWeight_1_weightRead_2_data[1639 : 1632];
  assign dSP_365_d = loadWeight_1_weightRead_2_data[1767 : 1760];
  assign dSP_365_b = _zz_b_2[103 : 96];
  assign dSP_366_a = loadWeight_1_weightRead_2_data[1647 : 1640];
  assign dSP_366_d = loadWeight_1_weightRead_2_data[1775 : 1768];
  assign dSP_366_b = _zz_b_2[111 : 104];
  assign dSP_367_a = loadWeight_1_weightRead_2_data[1655 : 1648];
  assign dSP_367_d = loadWeight_1_weightRead_2_data[1783 : 1776];
  assign dSP_367_b = _zz_b_2[119 : 112];
  assign dSP_368_a = loadWeight_1_weightRead_2_data[1663 : 1656];
  assign dSP_368_d = loadWeight_1_weightRead_2_data[1791 : 1784];
  assign dSP_368_b = _zz_b_2[127 : 120];
  assign dSP_369_a = loadWeight_1_weightRead_2_data[1799 : 1792];
  assign dSP_369_d = loadWeight_1_weightRead_2_data[1927 : 1920];
  assign dSP_369_b = _zz_b_2[7 : 0];
  assign dSP_370_a = loadWeight_1_weightRead_2_data[1807 : 1800];
  assign dSP_370_d = loadWeight_1_weightRead_2_data[1935 : 1928];
  assign dSP_370_b = _zz_b_2[15 : 8];
  assign dSP_371_a = loadWeight_1_weightRead_2_data[1815 : 1808];
  assign dSP_371_d = loadWeight_1_weightRead_2_data[1943 : 1936];
  assign dSP_371_b = _zz_b_2[23 : 16];
  assign dSP_372_a = loadWeight_1_weightRead_2_data[1823 : 1816];
  assign dSP_372_d = loadWeight_1_weightRead_2_data[1951 : 1944];
  assign dSP_372_b = _zz_b_2[31 : 24];
  assign dSP_373_a = loadWeight_1_weightRead_2_data[1831 : 1824];
  assign dSP_373_d = loadWeight_1_weightRead_2_data[1959 : 1952];
  assign dSP_373_b = _zz_b_2[39 : 32];
  assign dSP_374_a = loadWeight_1_weightRead_2_data[1839 : 1832];
  assign dSP_374_d = loadWeight_1_weightRead_2_data[1967 : 1960];
  assign dSP_374_b = _zz_b_2[47 : 40];
  assign dSP_375_a = loadWeight_1_weightRead_2_data[1847 : 1840];
  assign dSP_375_d = loadWeight_1_weightRead_2_data[1975 : 1968];
  assign dSP_375_b = _zz_b_2[55 : 48];
  assign dSP_376_a = loadWeight_1_weightRead_2_data[1855 : 1848];
  assign dSP_376_d = loadWeight_1_weightRead_2_data[1983 : 1976];
  assign dSP_376_b = _zz_b_2[63 : 56];
  assign dSP_377_a = loadWeight_1_weightRead_2_data[1863 : 1856];
  assign dSP_377_d = loadWeight_1_weightRead_2_data[1991 : 1984];
  assign dSP_377_b = _zz_b_2[71 : 64];
  assign dSP_378_a = loadWeight_1_weightRead_2_data[1871 : 1864];
  assign dSP_378_d = loadWeight_1_weightRead_2_data[1999 : 1992];
  assign dSP_378_b = _zz_b_2[79 : 72];
  assign dSP_379_a = loadWeight_1_weightRead_2_data[1879 : 1872];
  assign dSP_379_d = loadWeight_1_weightRead_2_data[2007 : 2000];
  assign dSP_379_b = _zz_b_2[87 : 80];
  assign dSP_380_a = loadWeight_1_weightRead_2_data[1887 : 1880];
  assign dSP_380_d = loadWeight_1_weightRead_2_data[2015 : 2008];
  assign dSP_380_b = _zz_b_2[95 : 88];
  assign dSP_381_a = loadWeight_1_weightRead_2_data[1895 : 1888];
  assign dSP_381_d = loadWeight_1_weightRead_2_data[2023 : 2016];
  assign dSP_381_b = _zz_b_2[103 : 96];
  assign dSP_382_a = loadWeight_1_weightRead_2_data[1903 : 1896];
  assign dSP_382_d = loadWeight_1_weightRead_2_data[2031 : 2024];
  assign dSP_382_b = _zz_b_2[111 : 104];
  assign dSP_383_a = loadWeight_1_weightRead_2_data[1911 : 1904];
  assign dSP_383_d = loadWeight_1_weightRead_2_data[2039 : 2032];
  assign dSP_383_b = _zz_b_2[119 : 112];
  assign dSP_384_a = loadWeight_1_weightRead_2_data[1919 : 1912];
  assign dSP_384_d = loadWeight_1_weightRead_2_data[2047 : 2040];
  assign dSP_384_b = _zz_b_2[127 : 120];
  assign dSP_385_a = loadWeight_1_weightRead_3_data[7 : 0];
  assign dSP_385_d = loadWeight_1_weightRead_3_data[135 : 128];
  assign dSP_385_b = _zz_b_3[7 : 0];
  assign dSP_386_a = loadWeight_1_weightRead_3_data[15 : 8];
  assign dSP_386_d = loadWeight_1_weightRead_3_data[143 : 136];
  assign dSP_386_b = _zz_b_3[15 : 8];
  assign dSP_387_a = loadWeight_1_weightRead_3_data[23 : 16];
  assign dSP_387_d = loadWeight_1_weightRead_3_data[151 : 144];
  assign dSP_387_b = _zz_b_3[23 : 16];
  assign dSP_388_a = loadWeight_1_weightRead_3_data[31 : 24];
  assign dSP_388_d = loadWeight_1_weightRead_3_data[159 : 152];
  assign dSP_388_b = _zz_b_3[31 : 24];
  assign dSP_389_a = loadWeight_1_weightRead_3_data[39 : 32];
  assign dSP_389_d = loadWeight_1_weightRead_3_data[167 : 160];
  assign dSP_389_b = _zz_b_3[39 : 32];
  assign dSP_390_a = loadWeight_1_weightRead_3_data[47 : 40];
  assign dSP_390_d = loadWeight_1_weightRead_3_data[175 : 168];
  assign dSP_390_b = _zz_b_3[47 : 40];
  assign dSP_391_a = loadWeight_1_weightRead_3_data[55 : 48];
  assign dSP_391_d = loadWeight_1_weightRead_3_data[183 : 176];
  assign dSP_391_b = _zz_b_3[55 : 48];
  assign dSP_392_a = loadWeight_1_weightRead_3_data[63 : 56];
  assign dSP_392_d = loadWeight_1_weightRead_3_data[191 : 184];
  assign dSP_392_b = _zz_b_3[63 : 56];
  assign dSP_393_a = loadWeight_1_weightRead_3_data[71 : 64];
  assign dSP_393_d = loadWeight_1_weightRead_3_data[199 : 192];
  assign dSP_393_b = _zz_b_3[71 : 64];
  assign dSP_394_a = loadWeight_1_weightRead_3_data[79 : 72];
  assign dSP_394_d = loadWeight_1_weightRead_3_data[207 : 200];
  assign dSP_394_b = _zz_b_3[79 : 72];
  assign dSP_395_a = loadWeight_1_weightRead_3_data[87 : 80];
  assign dSP_395_d = loadWeight_1_weightRead_3_data[215 : 208];
  assign dSP_395_b = _zz_b_3[87 : 80];
  assign dSP_396_a = loadWeight_1_weightRead_3_data[95 : 88];
  assign dSP_396_d = loadWeight_1_weightRead_3_data[223 : 216];
  assign dSP_396_b = _zz_b_3[95 : 88];
  assign dSP_397_a = loadWeight_1_weightRead_3_data[103 : 96];
  assign dSP_397_d = loadWeight_1_weightRead_3_data[231 : 224];
  assign dSP_397_b = _zz_b_3[103 : 96];
  assign dSP_398_a = loadWeight_1_weightRead_3_data[111 : 104];
  assign dSP_398_d = loadWeight_1_weightRead_3_data[239 : 232];
  assign dSP_398_b = _zz_b_3[111 : 104];
  assign dSP_399_a = loadWeight_1_weightRead_3_data[119 : 112];
  assign dSP_399_d = loadWeight_1_weightRead_3_data[247 : 240];
  assign dSP_399_b = _zz_b_3[119 : 112];
  assign dSP_400_a = loadWeight_1_weightRead_3_data[127 : 120];
  assign dSP_400_d = loadWeight_1_weightRead_3_data[255 : 248];
  assign dSP_400_b = _zz_b_3[127 : 120];
  assign dSP_401_a = loadWeight_1_weightRead_3_data[263 : 256];
  assign dSP_401_d = loadWeight_1_weightRead_3_data[391 : 384];
  assign dSP_401_b = _zz_b_3[7 : 0];
  assign dSP_402_a = loadWeight_1_weightRead_3_data[271 : 264];
  assign dSP_402_d = loadWeight_1_weightRead_3_data[399 : 392];
  assign dSP_402_b = _zz_b_3[15 : 8];
  assign dSP_403_a = loadWeight_1_weightRead_3_data[279 : 272];
  assign dSP_403_d = loadWeight_1_weightRead_3_data[407 : 400];
  assign dSP_403_b = _zz_b_3[23 : 16];
  assign dSP_404_a = loadWeight_1_weightRead_3_data[287 : 280];
  assign dSP_404_d = loadWeight_1_weightRead_3_data[415 : 408];
  assign dSP_404_b = _zz_b_3[31 : 24];
  assign dSP_405_a = loadWeight_1_weightRead_3_data[295 : 288];
  assign dSP_405_d = loadWeight_1_weightRead_3_data[423 : 416];
  assign dSP_405_b = _zz_b_3[39 : 32];
  assign dSP_406_a = loadWeight_1_weightRead_3_data[303 : 296];
  assign dSP_406_d = loadWeight_1_weightRead_3_data[431 : 424];
  assign dSP_406_b = _zz_b_3[47 : 40];
  assign dSP_407_a = loadWeight_1_weightRead_3_data[311 : 304];
  assign dSP_407_d = loadWeight_1_weightRead_3_data[439 : 432];
  assign dSP_407_b = _zz_b_3[55 : 48];
  assign dSP_408_a = loadWeight_1_weightRead_3_data[319 : 312];
  assign dSP_408_d = loadWeight_1_weightRead_3_data[447 : 440];
  assign dSP_408_b = _zz_b_3[63 : 56];
  assign dSP_409_a = loadWeight_1_weightRead_3_data[327 : 320];
  assign dSP_409_d = loadWeight_1_weightRead_3_data[455 : 448];
  assign dSP_409_b = _zz_b_3[71 : 64];
  assign dSP_410_a = loadWeight_1_weightRead_3_data[335 : 328];
  assign dSP_410_d = loadWeight_1_weightRead_3_data[463 : 456];
  assign dSP_410_b = _zz_b_3[79 : 72];
  assign dSP_411_a = loadWeight_1_weightRead_3_data[343 : 336];
  assign dSP_411_d = loadWeight_1_weightRead_3_data[471 : 464];
  assign dSP_411_b = _zz_b_3[87 : 80];
  assign dSP_412_a = loadWeight_1_weightRead_3_data[351 : 344];
  assign dSP_412_d = loadWeight_1_weightRead_3_data[479 : 472];
  assign dSP_412_b = _zz_b_3[95 : 88];
  assign dSP_413_a = loadWeight_1_weightRead_3_data[359 : 352];
  assign dSP_413_d = loadWeight_1_weightRead_3_data[487 : 480];
  assign dSP_413_b = _zz_b_3[103 : 96];
  assign dSP_414_a = loadWeight_1_weightRead_3_data[367 : 360];
  assign dSP_414_d = loadWeight_1_weightRead_3_data[495 : 488];
  assign dSP_414_b = _zz_b_3[111 : 104];
  assign dSP_415_a = loadWeight_1_weightRead_3_data[375 : 368];
  assign dSP_415_d = loadWeight_1_weightRead_3_data[503 : 496];
  assign dSP_415_b = _zz_b_3[119 : 112];
  assign dSP_416_a = loadWeight_1_weightRead_3_data[383 : 376];
  assign dSP_416_d = loadWeight_1_weightRead_3_data[511 : 504];
  assign dSP_416_b = _zz_b_3[127 : 120];
  assign dSP_417_a = loadWeight_1_weightRead_3_data[519 : 512];
  assign dSP_417_d = loadWeight_1_weightRead_3_data[647 : 640];
  assign dSP_417_b = _zz_b_3[7 : 0];
  assign dSP_418_a = loadWeight_1_weightRead_3_data[527 : 520];
  assign dSP_418_d = loadWeight_1_weightRead_3_data[655 : 648];
  assign dSP_418_b = _zz_b_3[15 : 8];
  assign dSP_419_a = loadWeight_1_weightRead_3_data[535 : 528];
  assign dSP_419_d = loadWeight_1_weightRead_3_data[663 : 656];
  assign dSP_419_b = _zz_b_3[23 : 16];
  assign dSP_420_a = loadWeight_1_weightRead_3_data[543 : 536];
  assign dSP_420_d = loadWeight_1_weightRead_3_data[671 : 664];
  assign dSP_420_b = _zz_b_3[31 : 24];
  assign dSP_421_a = loadWeight_1_weightRead_3_data[551 : 544];
  assign dSP_421_d = loadWeight_1_weightRead_3_data[679 : 672];
  assign dSP_421_b = _zz_b_3[39 : 32];
  assign dSP_422_a = loadWeight_1_weightRead_3_data[559 : 552];
  assign dSP_422_d = loadWeight_1_weightRead_3_data[687 : 680];
  assign dSP_422_b = _zz_b_3[47 : 40];
  assign dSP_423_a = loadWeight_1_weightRead_3_data[567 : 560];
  assign dSP_423_d = loadWeight_1_weightRead_3_data[695 : 688];
  assign dSP_423_b = _zz_b_3[55 : 48];
  assign dSP_424_a = loadWeight_1_weightRead_3_data[575 : 568];
  assign dSP_424_d = loadWeight_1_weightRead_3_data[703 : 696];
  assign dSP_424_b = _zz_b_3[63 : 56];
  assign dSP_425_a = loadWeight_1_weightRead_3_data[583 : 576];
  assign dSP_425_d = loadWeight_1_weightRead_3_data[711 : 704];
  assign dSP_425_b = _zz_b_3[71 : 64];
  assign dSP_426_a = loadWeight_1_weightRead_3_data[591 : 584];
  assign dSP_426_d = loadWeight_1_weightRead_3_data[719 : 712];
  assign dSP_426_b = _zz_b_3[79 : 72];
  assign dSP_427_a = loadWeight_1_weightRead_3_data[599 : 592];
  assign dSP_427_d = loadWeight_1_weightRead_3_data[727 : 720];
  assign dSP_427_b = _zz_b_3[87 : 80];
  assign dSP_428_a = loadWeight_1_weightRead_3_data[607 : 600];
  assign dSP_428_d = loadWeight_1_weightRead_3_data[735 : 728];
  assign dSP_428_b = _zz_b_3[95 : 88];
  assign dSP_429_a = loadWeight_1_weightRead_3_data[615 : 608];
  assign dSP_429_d = loadWeight_1_weightRead_3_data[743 : 736];
  assign dSP_429_b = _zz_b_3[103 : 96];
  assign dSP_430_a = loadWeight_1_weightRead_3_data[623 : 616];
  assign dSP_430_d = loadWeight_1_weightRead_3_data[751 : 744];
  assign dSP_430_b = _zz_b_3[111 : 104];
  assign dSP_431_a = loadWeight_1_weightRead_3_data[631 : 624];
  assign dSP_431_d = loadWeight_1_weightRead_3_data[759 : 752];
  assign dSP_431_b = _zz_b_3[119 : 112];
  assign dSP_432_a = loadWeight_1_weightRead_3_data[639 : 632];
  assign dSP_432_d = loadWeight_1_weightRead_3_data[767 : 760];
  assign dSP_432_b = _zz_b_3[127 : 120];
  assign dSP_433_a = loadWeight_1_weightRead_3_data[775 : 768];
  assign dSP_433_d = loadWeight_1_weightRead_3_data[903 : 896];
  assign dSP_433_b = _zz_b_3[7 : 0];
  assign dSP_434_a = loadWeight_1_weightRead_3_data[783 : 776];
  assign dSP_434_d = loadWeight_1_weightRead_3_data[911 : 904];
  assign dSP_434_b = _zz_b_3[15 : 8];
  assign dSP_435_a = loadWeight_1_weightRead_3_data[791 : 784];
  assign dSP_435_d = loadWeight_1_weightRead_3_data[919 : 912];
  assign dSP_435_b = _zz_b_3[23 : 16];
  assign dSP_436_a = loadWeight_1_weightRead_3_data[799 : 792];
  assign dSP_436_d = loadWeight_1_weightRead_3_data[927 : 920];
  assign dSP_436_b = _zz_b_3[31 : 24];
  assign dSP_437_a = loadWeight_1_weightRead_3_data[807 : 800];
  assign dSP_437_d = loadWeight_1_weightRead_3_data[935 : 928];
  assign dSP_437_b = _zz_b_3[39 : 32];
  assign dSP_438_a = loadWeight_1_weightRead_3_data[815 : 808];
  assign dSP_438_d = loadWeight_1_weightRead_3_data[943 : 936];
  assign dSP_438_b = _zz_b_3[47 : 40];
  assign dSP_439_a = loadWeight_1_weightRead_3_data[823 : 816];
  assign dSP_439_d = loadWeight_1_weightRead_3_data[951 : 944];
  assign dSP_439_b = _zz_b_3[55 : 48];
  assign dSP_440_a = loadWeight_1_weightRead_3_data[831 : 824];
  assign dSP_440_d = loadWeight_1_weightRead_3_data[959 : 952];
  assign dSP_440_b = _zz_b_3[63 : 56];
  assign dSP_441_a = loadWeight_1_weightRead_3_data[839 : 832];
  assign dSP_441_d = loadWeight_1_weightRead_3_data[967 : 960];
  assign dSP_441_b = _zz_b_3[71 : 64];
  assign dSP_442_a = loadWeight_1_weightRead_3_data[847 : 840];
  assign dSP_442_d = loadWeight_1_weightRead_3_data[975 : 968];
  assign dSP_442_b = _zz_b_3[79 : 72];
  assign dSP_443_a = loadWeight_1_weightRead_3_data[855 : 848];
  assign dSP_443_d = loadWeight_1_weightRead_3_data[983 : 976];
  assign dSP_443_b = _zz_b_3[87 : 80];
  assign dSP_444_a = loadWeight_1_weightRead_3_data[863 : 856];
  assign dSP_444_d = loadWeight_1_weightRead_3_data[991 : 984];
  assign dSP_444_b = _zz_b_3[95 : 88];
  assign dSP_445_a = loadWeight_1_weightRead_3_data[871 : 864];
  assign dSP_445_d = loadWeight_1_weightRead_3_data[999 : 992];
  assign dSP_445_b = _zz_b_3[103 : 96];
  assign dSP_446_a = loadWeight_1_weightRead_3_data[879 : 872];
  assign dSP_446_d = loadWeight_1_weightRead_3_data[1007 : 1000];
  assign dSP_446_b = _zz_b_3[111 : 104];
  assign dSP_447_a = loadWeight_1_weightRead_3_data[887 : 880];
  assign dSP_447_d = loadWeight_1_weightRead_3_data[1015 : 1008];
  assign dSP_447_b = _zz_b_3[119 : 112];
  assign dSP_448_a = loadWeight_1_weightRead_3_data[895 : 888];
  assign dSP_448_d = loadWeight_1_weightRead_3_data[1023 : 1016];
  assign dSP_448_b = _zz_b_3[127 : 120];
  assign dSP_449_a = loadWeight_1_weightRead_3_data[1031 : 1024];
  assign dSP_449_d = loadWeight_1_weightRead_3_data[1159 : 1152];
  assign dSP_449_b = _zz_b_3[7 : 0];
  assign dSP_450_a = loadWeight_1_weightRead_3_data[1039 : 1032];
  assign dSP_450_d = loadWeight_1_weightRead_3_data[1167 : 1160];
  assign dSP_450_b = _zz_b_3[15 : 8];
  assign dSP_451_a = loadWeight_1_weightRead_3_data[1047 : 1040];
  assign dSP_451_d = loadWeight_1_weightRead_3_data[1175 : 1168];
  assign dSP_451_b = _zz_b_3[23 : 16];
  assign dSP_452_a = loadWeight_1_weightRead_3_data[1055 : 1048];
  assign dSP_452_d = loadWeight_1_weightRead_3_data[1183 : 1176];
  assign dSP_452_b = _zz_b_3[31 : 24];
  assign dSP_453_a = loadWeight_1_weightRead_3_data[1063 : 1056];
  assign dSP_453_d = loadWeight_1_weightRead_3_data[1191 : 1184];
  assign dSP_453_b = _zz_b_3[39 : 32];
  assign dSP_454_a = loadWeight_1_weightRead_3_data[1071 : 1064];
  assign dSP_454_d = loadWeight_1_weightRead_3_data[1199 : 1192];
  assign dSP_454_b = _zz_b_3[47 : 40];
  assign dSP_455_a = loadWeight_1_weightRead_3_data[1079 : 1072];
  assign dSP_455_d = loadWeight_1_weightRead_3_data[1207 : 1200];
  assign dSP_455_b = _zz_b_3[55 : 48];
  assign dSP_456_a = loadWeight_1_weightRead_3_data[1087 : 1080];
  assign dSP_456_d = loadWeight_1_weightRead_3_data[1215 : 1208];
  assign dSP_456_b = _zz_b_3[63 : 56];
  assign dSP_457_a = loadWeight_1_weightRead_3_data[1095 : 1088];
  assign dSP_457_d = loadWeight_1_weightRead_3_data[1223 : 1216];
  assign dSP_457_b = _zz_b_3[71 : 64];
  assign dSP_458_a = loadWeight_1_weightRead_3_data[1103 : 1096];
  assign dSP_458_d = loadWeight_1_weightRead_3_data[1231 : 1224];
  assign dSP_458_b = _zz_b_3[79 : 72];
  assign dSP_459_a = loadWeight_1_weightRead_3_data[1111 : 1104];
  assign dSP_459_d = loadWeight_1_weightRead_3_data[1239 : 1232];
  assign dSP_459_b = _zz_b_3[87 : 80];
  assign dSP_460_a = loadWeight_1_weightRead_3_data[1119 : 1112];
  assign dSP_460_d = loadWeight_1_weightRead_3_data[1247 : 1240];
  assign dSP_460_b = _zz_b_3[95 : 88];
  assign dSP_461_a = loadWeight_1_weightRead_3_data[1127 : 1120];
  assign dSP_461_d = loadWeight_1_weightRead_3_data[1255 : 1248];
  assign dSP_461_b = _zz_b_3[103 : 96];
  assign dSP_462_a = loadWeight_1_weightRead_3_data[1135 : 1128];
  assign dSP_462_d = loadWeight_1_weightRead_3_data[1263 : 1256];
  assign dSP_462_b = _zz_b_3[111 : 104];
  assign dSP_463_a = loadWeight_1_weightRead_3_data[1143 : 1136];
  assign dSP_463_d = loadWeight_1_weightRead_3_data[1271 : 1264];
  assign dSP_463_b = _zz_b_3[119 : 112];
  assign dSP_464_a = loadWeight_1_weightRead_3_data[1151 : 1144];
  assign dSP_464_d = loadWeight_1_weightRead_3_data[1279 : 1272];
  assign dSP_464_b = _zz_b_3[127 : 120];
  assign dSP_465_a = loadWeight_1_weightRead_3_data[1287 : 1280];
  assign dSP_465_d = loadWeight_1_weightRead_3_data[1415 : 1408];
  assign dSP_465_b = _zz_b_3[7 : 0];
  assign dSP_466_a = loadWeight_1_weightRead_3_data[1295 : 1288];
  assign dSP_466_d = loadWeight_1_weightRead_3_data[1423 : 1416];
  assign dSP_466_b = _zz_b_3[15 : 8];
  assign dSP_467_a = loadWeight_1_weightRead_3_data[1303 : 1296];
  assign dSP_467_d = loadWeight_1_weightRead_3_data[1431 : 1424];
  assign dSP_467_b = _zz_b_3[23 : 16];
  assign dSP_468_a = loadWeight_1_weightRead_3_data[1311 : 1304];
  assign dSP_468_d = loadWeight_1_weightRead_3_data[1439 : 1432];
  assign dSP_468_b = _zz_b_3[31 : 24];
  assign dSP_469_a = loadWeight_1_weightRead_3_data[1319 : 1312];
  assign dSP_469_d = loadWeight_1_weightRead_3_data[1447 : 1440];
  assign dSP_469_b = _zz_b_3[39 : 32];
  assign dSP_470_a = loadWeight_1_weightRead_3_data[1327 : 1320];
  assign dSP_470_d = loadWeight_1_weightRead_3_data[1455 : 1448];
  assign dSP_470_b = _zz_b_3[47 : 40];
  assign dSP_471_a = loadWeight_1_weightRead_3_data[1335 : 1328];
  assign dSP_471_d = loadWeight_1_weightRead_3_data[1463 : 1456];
  assign dSP_471_b = _zz_b_3[55 : 48];
  assign dSP_472_a = loadWeight_1_weightRead_3_data[1343 : 1336];
  assign dSP_472_d = loadWeight_1_weightRead_3_data[1471 : 1464];
  assign dSP_472_b = _zz_b_3[63 : 56];
  assign dSP_473_a = loadWeight_1_weightRead_3_data[1351 : 1344];
  assign dSP_473_d = loadWeight_1_weightRead_3_data[1479 : 1472];
  assign dSP_473_b = _zz_b_3[71 : 64];
  assign dSP_474_a = loadWeight_1_weightRead_3_data[1359 : 1352];
  assign dSP_474_d = loadWeight_1_weightRead_3_data[1487 : 1480];
  assign dSP_474_b = _zz_b_3[79 : 72];
  assign dSP_475_a = loadWeight_1_weightRead_3_data[1367 : 1360];
  assign dSP_475_d = loadWeight_1_weightRead_3_data[1495 : 1488];
  assign dSP_475_b = _zz_b_3[87 : 80];
  assign dSP_476_a = loadWeight_1_weightRead_3_data[1375 : 1368];
  assign dSP_476_d = loadWeight_1_weightRead_3_data[1503 : 1496];
  assign dSP_476_b = _zz_b_3[95 : 88];
  assign dSP_477_a = loadWeight_1_weightRead_3_data[1383 : 1376];
  assign dSP_477_d = loadWeight_1_weightRead_3_data[1511 : 1504];
  assign dSP_477_b = _zz_b_3[103 : 96];
  assign dSP_478_a = loadWeight_1_weightRead_3_data[1391 : 1384];
  assign dSP_478_d = loadWeight_1_weightRead_3_data[1519 : 1512];
  assign dSP_478_b = _zz_b_3[111 : 104];
  assign dSP_479_a = loadWeight_1_weightRead_3_data[1399 : 1392];
  assign dSP_479_d = loadWeight_1_weightRead_3_data[1527 : 1520];
  assign dSP_479_b = _zz_b_3[119 : 112];
  assign dSP_480_a = loadWeight_1_weightRead_3_data[1407 : 1400];
  assign dSP_480_d = loadWeight_1_weightRead_3_data[1535 : 1528];
  assign dSP_480_b = _zz_b_3[127 : 120];
  assign dSP_481_a = loadWeight_1_weightRead_3_data[1543 : 1536];
  assign dSP_481_d = loadWeight_1_weightRead_3_data[1671 : 1664];
  assign dSP_481_b = _zz_b_3[7 : 0];
  assign dSP_482_a = loadWeight_1_weightRead_3_data[1551 : 1544];
  assign dSP_482_d = loadWeight_1_weightRead_3_data[1679 : 1672];
  assign dSP_482_b = _zz_b_3[15 : 8];
  assign dSP_483_a = loadWeight_1_weightRead_3_data[1559 : 1552];
  assign dSP_483_d = loadWeight_1_weightRead_3_data[1687 : 1680];
  assign dSP_483_b = _zz_b_3[23 : 16];
  assign dSP_484_a = loadWeight_1_weightRead_3_data[1567 : 1560];
  assign dSP_484_d = loadWeight_1_weightRead_3_data[1695 : 1688];
  assign dSP_484_b = _zz_b_3[31 : 24];
  assign dSP_485_a = loadWeight_1_weightRead_3_data[1575 : 1568];
  assign dSP_485_d = loadWeight_1_weightRead_3_data[1703 : 1696];
  assign dSP_485_b = _zz_b_3[39 : 32];
  assign dSP_486_a = loadWeight_1_weightRead_3_data[1583 : 1576];
  assign dSP_486_d = loadWeight_1_weightRead_3_data[1711 : 1704];
  assign dSP_486_b = _zz_b_3[47 : 40];
  assign dSP_487_a = loadWeight_1_weightRead_3_data[1591 : 1584];
  assign dSP_487_d = loadWeight_1_weightRead_3_data[1719 : 1712];
  assign dSP_487_b = _zz_b_3[55 : 48];
  assign dSP_488_a = loadWeight_1_weightRead_3_data[1599 : 1592];
  assign dSP_488_d = loadWeight_1_weightRead_3_data[1727 : 1720];
  assign dSP_488_b = _zz_b_3[63 : 56];
  assign dSP_489_a = loadWeight_1_weightRead_3_data[1607 : 1600];
  assign dSP_489_d = loadWeight_1_weightRead_3_data[1735 : 1728];
  assign dSP_489_b = _zz_b_3[71 : 64];
  assign dSP_490_a = loadWeight_1_weightRead_3_data[1615 : 1608];
  assign dSP_490_d = loadWeight_1_weightRead_3_data[1743 : 1736];
  assign dSP_490_b = _zz_b_3[79 : 72];
  assign dSP_491_a = loadWeight_1_weightRead_3_data[1623 : 1616];
  assign dSP_491_d = loadWeight_1_weightRead_3_data[1751 : 1744];
  assign dSP_491_b = _zz_b_3[87 : 80];
  assign dSP_492_a = loadWeight_1_weightRead_3_data[1631 : 1624];
  assign dSP_492_d = loadWeight_1_weightRead_3_data[1759 : 1752];
  assign dSP_492_b = _zz_b_3[95 : 88];
  assign dSP_493_a = loadWeight_1_weightRead_3_data[1639 : 1632];
  assign dSP_493_d = loadWeight_1_weightRead_3_data[1767 : 1760];
  assign dSP_493_b = _zz_b_3[103 : 96];
  assign dSP_494_a = loadWeight_1_weightRead_3_data[1647 : 1640];
  assign dSP_494_d = loadWeight_1_weightRead_3_data[1775 : 1768];
  assign dSP_494_b = _zz_b_3[111 : 104];
  assign dSP_495_a = loadWeight_1_weightRead_3_data[1655 : 1648];
  assign dSP_495_d = loadWeight_1_weightRead_3_data[1783 : 1776];
  assign dSP_495_b = _zz_b_3[119 : 112];
  assign dSP_496_a = loadWeight_1_weightRead_3_data[1663 : 1656];
  assign dSP_496_d = loadWeight_1_weightRead_3_data[1791 : 1784];
  assign dSP_496_b = _zz_b_3[127 : 120];
  assign dSP_497_a = loadWeight_1_weightRead_3_data[1799 : 1792];
  assign dSP_497_d = loadWeight_1_weightRead_3_data[1927 : 1920];
  assign dSP_497_b = _zz_b_3[7 : 0];
  assign dSP_498_a = loadWeight_1_weightRead_3_data[1807 : 1800];
  assign dSP_498_d = loadWeight_1_weightRead_3_data[1935 : 1928];
  assign dSP_498_b = _zz_b_3[15 : 8];
  assign dSP_499_a = loadWeight_1_weightRead_3_data[1815 : 1808];
  assign dSP_499_d = loadWeight_1_weightRead_3_data[1943 : 1936];
  assign dSP_499_b = _zz_b_3[23 : 16];
  assign dSP_500_a = loadWeight_1_weightRead_3_data[1823 : 1816];
  assign dSP_500_d = loadWeight_1_weightRead_3_data[1951 : 1944];
  assign dSP_500_b = _zz_b_3[31 : 24];
  assign dSP_501_a = loadWeight_1_weightRead_3_data[1831 : 1824];
  assign dSP_501_d = loadWeight_1_weightRead_3_data[1959 : 1952];
  assign dSP_501_b = _zz_b_3[39 : 32];
  assign dSP_502_a = loadWeight_1_weightRead_3_data[1839 : 1832];
  assign dSP_502_d = loadWeight_1_weightRead_3_data[1967 : 1960];
  assign dSP_502_b = _zz_b_3[47 : 40];
  assign dSP_503_a = loadWeight_1_weightRead_3_data[1847 : 1840];
  assign dSP_503_d = loadWeight_1_weightRead_3_data[1975 : 1968];
  assign dSP_503_b = _zz_b_3[55 : 48];
  assign dSP_504_a = loadWeight_1_weightRead_3_data[1855 : 1848];
  assign dSP_504_d = loadWeight_1_weightRead_3_data[1983 : 1976];
  assign dSP_504_b = _zz_b_3[63 : 56];
  assign dSP_505_a = loadWeight_1_weightRead_3_data[1863 : 1856];
  assign dSP_505_d = loadWeight_1_weightRead_3_data[1991 : 1984];
  assign dSP_505_b = _zz_b_3[71 : 64];
  assign dSP_506_a = loadWeight_1_weightRead_3_data[1871 : 1864];
  assign dSP_506_d = loadWeight_1_weightRead_3_data[1999 : 1992];
  assign dSP_506_b = _zz_b_3[79 : 72];
  assign dSP_507_a = loadWeight_1_weightRead_3_data[1879 : 1872];
  assign dSP_507_d = loadWeight_1_weightRead_3_data[2007 : 2000];
  assign dSP_507_b = _zz_b_3[87 : 80];
  assign dSP_508_a = loadWeight_1_weightRead_3_data[1887 : 1880];
  assign dSP_508_d = loadWeight_1_weightRead_3_data[2015 : 2008];
  assign dSP_508_b = _zz_b_3[95 : 88];
  assign dSP_509_a = loadWeight_1_weightRead_3_data[1895 : 1888];
  assign dSP_509_d = loadWeight_1_weightRead_3_data[2023 : 2016];
  assign dSP_509_b = _zz_b_3[103 : 96];
  assign dSP_510_a = loadWeight_1_weightRead_3_data[1903 : 1896];
  assign dSP_510_d = loadWeight_1_weightRead_3_data[2031 : 2024];
  assign dSP_510_b = _zz_b_3[111 : 104];
  assign dSP_511_a = loadWeight_1_weightRead_3_data[1911 : 1904];
  assign dSP_511_d = loadWeight_1_weightRead_3_data[2039 : 2032];
  assign dSP_511_b = _zz_b_3[119 : 112];
  assign dSP_512_a = loadWeight_1_weightRead_3_data[1919 : 1912];
  assign dSP_512_d = loadWeight_1_weightRead_3_data[2047 : 2040];
  assign dSP_512_b = _zz_b_3[127 : 120];
  assign dSP_513_a = loadWeight_1_weightRead_4_data[7 : 0];
  assign dSP_513_d = loadWeight_1_weightRead_4_data[135 : 128];
  assign dSP_513_b = _zz_b_4[7 : 0];
  assign dSP_514_a = loadWeight_1_weightRead_4_data[15 : 8];
  assign dSP_514_d = loadWeight_1_weightRead_4_data[143 : 136];
  assign dSP_514_b = _zz_b_4[15 : 8];
  assign dSP_515_a = loadWeight_1_weightRead_4_data[23 : 16];
  assign dSP_515_d = loadWeight_1_weightRead_4_data[151 : 144];
  assign dSP_515_b = _zz_b_4[23 : 16];
  assign dSP_516_a = loadWeight_1_weightRead_4_data[31 : 24];
  assign dSP_516_d = loadWeight_1_weightRead_4_data[159 : 152];
  assign dSP_516_b = _zz_b_4[31 : 24];
  assign dSP_517_a = loadWeight_1_weightRead_4_data[39 : 32];
  assign dSP_517_d = loadWeight_1_weightRead_4_data[167 : 160];
  assign dSP_517_b = _zz_b_4[39 : 32];
  assign dSP_518_a = loadWeight_1_weightRead_4_data[47 : 40];
  assign dSP_518_d = loadWeight_1_weightRead_4_data[175 : 168];
  assign dSP_518_b = _zz_b_4[47 : 40];
  assign dSP_519_a = loadWeight_1_weightRead_4_data[55 : 48];
  assign dSP_519_d = loadWeight_1_weightRead_4_data[183 : 176];
  assign dSP_519_b = _zz_b_4[55 : 48];
  assign dSP_520_a = loadWeight_1_weightRead_4_data[63 : 56];
  assign dSP_520_d = loadWeight_1_weightRead_4_data[191 : 184];
  assign dSP_520_b = _zz_b_4[63 : 56];
  assign dSP_521_a = loadWeight_1_weightRead_4_data[71 : 64];
  assign dSP_521_d = loadWeight_1_weightRead_4_data[199 : 192];
  assign dSP_521_b = _zz_b_4[71 : 64];
  assign dSP_522_a = loadWeight_1_weightRead_4_data[79 : 72];
  assign dSP_522_d = loadWeight_1_weightRead_4_data[207 : 200];
  assign dSP_522_b = _zz_b_4[79 : 72];
  assign dSP_523_a = loadWeight_1_weightRead_4_data[87 : 80];
  assign dSP_523_d = loadWeight_1_weightRead_4_data[215 : 208];
  assign dSP_523_b = _zz_b_4[87 : 80];
  assign dSP_524_a = loadWeight_1_weightRead_4_data[95 : 88];
  assign dSP_524_d = loadWeight_1_weightRead_4_data[223 : 216];
  assign dSP_524_b = _zz_b_4[95 : 88];
  assign dSP_525_a = loadWeight_1_weightRead_4_data[103 : 96];
  assign dSP_525_d = loadWeight_1_weightRead_4_data[231 : 224];
  assign dSP_525_b = _zz_b_4[103 : 96];
  assign dSP_526_a = loadWeight_1_weightRead_4_data[111 : 104];
  assign dSP_526_d = loadWeight_1_weightRead_4_data[239 : 232];
  assign dSP_526_b = _zz_b_4[111 : 104];
  assign dSP_527_a = loadWeight_1_weightRead_4_data[119 : 112];
  assign dSP_527_d = loadWeight_1_weightRead_4_data[247 : 240];
  assign dSP_527_b = _zz_b_4[119 : 112];
  assign dSP_528_a = loadWeight_1_weightRead_4_data[127 : 120];
  assign dSP_528_d = loadWeight_1_weightRead_4_data[255 : 248];
  assign dSP_528_b = _zz_b_4[127 : 120];
  assign dSP_529_a = loadWeight_1_weightRead_4_data[263 : 256];
  assign dSP_529_d = loadWeight_1_weightRead_4_data[391 : 384];
  assign dSP_529_b = _zz_b_4[7 : 0];
  assign dSP_530_a = loadWeight_1_weightRead_4_data[271 : 264];
  assign dSP_530_d = loadWeight_1_weightRead_4_data[399 : 392];
  assign dSP_530_b = _zz_b_4[15 : 8];
  assign dSP_531_a = loadWeight_1_weightRead_4_data[279 : 272];
  assign dSP_531_d = loadWeight_1_weightRead_4_data[407 : 400];
  assign dSP_531_b = _zz_b_4[23 : 16];
  assign dSP_532_a = loadWeight_1_weightRead_4_data[287 : 280];
  assign dSP_532_d = loadWeight_1_weightRead_4_data[415 : 408];
  assign dSP_532_b = _zz_b_4[31 : 24];
  assign dSP_533_a = loadWeight_1_weightRead_4_data[295 : 288];
  assign dSP_533_d = loadWeight_1_weightRead_4_data[423 : 416];
  assign dSP_533_b = _zz_b_4[39 : 32];
  assign dSP_534_a = loadWeight_1_weightRead_4_data[303 : 296];
  assign dSP_534_d = loadWeight_1_weightRead_4_data[431 : 424];
  assign dSP_534_b = _zz_b_4[47 : 40];
  assign dSP_535_a = loadWeight_1_weightRead_4_data[311 : 304];
  assign dSP_535_d = loadWeight_1_weightRead_4_data[439 : 432];
  assign dSP_535_b = _zz_b_4[55 : 48];
  assign dSP_536_a = loadWeight_1_weightRead_4_data[319 : 312];
  assign dSP_536_d = loadWeight_1_weightRead_4_data[447 : 440];
  assign dSP_536_b = _zz_b_4[63 : 56];
  assign dSP_537_a = loadWeight_1_weightRead_4_data[327 : 320];
  assign dSP_537_d = loadWeight_1_weightRead_4_data[455 : 448];
  assign dSP_537_b = _zz_b_4[71 : 64];
  assign dSP_538_a = loadWeight_1_weightRead_4_data[335 : 328];
  assign dSP_538_d = loadWeight_1_weightRead_4_data[463 : 456];
  assign dSP_538_b = _zz_b_4[79 : 72];
  assign dSP_539_a = loadWeight_1_weightRead_4_data[343 : 336];
  assign dSP_539_d = loadWeight_1_weightRead_4_data[471 : 464];
  assign dSP_539_b = _zz_b_4[87 : 80];
  assign dSP_540_a = loadWeight_1_weightRead_4_data[351 : 344];
  assign dSP_540_d = loadWeight_1_weightRead_4_data[479 : 472];
  assign dSP_540_b = _zz_b_4[95 : 88];
  assign dSP_541_a = loadWeight_1_weightRead_4_data[359 : 352];
  assign dSP_541_d = loadWeight_1_weightRead_4_data[487 : 480];
  assign dSP_541_b = _zz_b_4[103 : 96];
  assign dSP_542_a = loadWeight_1_weightRead_4_data[367 : 360];
  assign dSP_542_d = loadWeight_1_weightRead_4_data[495 : 488];
  assign dSP_542_b = _zz_b_4[111 : 104];
  assign dSP_543_a = loadWeight_1_weightRead_4_data[375 : 368];
  assign dSP_543_d = loadWeight_1_weightRead_4_data[503 : 496];
  assign dSP_543_b = _zz_b_4[119 : 112];
  assign dSP_544_a = loadWeight_1_weightRead_4_data[383 : 376];
  assign dSP_544_d = loadWeight_1_weightRead_4_data[511 : 504];
  assign dSP_544_b = _zz_b_4[127 : 120];
  assign dSP_545_a = loadWeight_1_weightRead_4_data[519 : 512];
  assign dSP_545_d = loadWeight_1_weightRead_4_data[647 : 640];
  assign dSP_545_b = _zz_b_4[7 : 0];
  assign dSP_546_a = loadWeight_1_weightRead_4_data[527 : 520];
  assign dSP_546_d = loadWeight_1_weightRead_4_data[655 : 648];
  assign dSP_546_b = _zz_b_4[15 : 8];
  assign dSP_547_a = loadWeight_1_weightRead_4_data[535 : 528];
  assign dSP_547_d = loadWeight_1_weightRead_4_data[663 : 656];
  assign dSP_547_b = _zz_b_4[23 : 16];
  assign dSP_548_a = loadWeight_1_weightRead_4_data[543 : 536];
  assign dSP_548_d = loadWeight_1_weightRead_4_data[671 : 664];
  assign dSP_548_b = _zz_b_4[31 : 24];
  assign dSP_549_a = loadWeight_1_weightRead_4_data[551 : 544];
  assign dSP_549_d = loadWeight_1_weightRead_4_data[679 : 672];
  assign dSP_549_b = _zz_b_4[39 : 32];
  assign dSP_550_a = loadWeight_1_weightRead_4_data[559 : 552];
  assign dSP_550_d = loadWeight_1_weightRead_4_data[687 : 680];
  assign dSP_550_b = _zz_b_4[47 : 40];
  assign dSP_551_a = loadWeight_1_weightRead_4_data[567 : 560];
  assign dSP_551_d = loadWeight_1_weightRead_4_data[695 : 688];
  assign dSP_551_b = _zz_b_4[55 : 48];
  assign dSP_552_a = loadWeight_1_weightRead_4_data[575 : 568];
  assign dSP_552_d = loadWeight_1_weightRead_4_data[703 : 696];
  assign dSP_552_b = _zz_b_4[63 : 56];
  assign dSP_553_a = loadWeight_1_weightRead_4_data[583 : 576];
  assign dSP_553_d = loadWeight_1_weightRead_4_data[711 : 704];
  assign dSP_553_b = _zz_b_4[71 : 64];
  assign dSP_554_a = loadWeight_1_weightRead_4_data[591 : 584];
  assign dSP_554_d = loadWeight_1_weightRead_4_data[719 : 712];
  assign dSP_554_b = _zz_b_4[79 : 72];
  assign dSP_555_a = loadWeight_1_weightRead_4_data[599 : 592];
  assign dSP_555_d = loadWeight_1_weightRead_4_data[727 : 720];
  assign dSP_555_b = _zz_b_4[87 : 80];
  assign dSP_556_a = loadWeight_1_weightRead_4_data[607 : 600];
  assign dSP_556_d = loadWeight_1_weightRead_4_data[735 : 728];
  assign dSP_556_b = _zz_b_4[95 : 88];
  assign dSP_557_a = loadWeight_1_weightRead_4_data[615 : 608];
  assign dSP_557_d = loadWeight_1_weightRead_4_data[743 : 736];
  assign dSP_557_b = _zz_b_4[103 : 96];
  assign dSP_558_a = loadWeight_1_weightRead_4_data[623 : 616];
  assign dSP_558_d = loadWeight_1_weightRead_4_data[751 : 744];
  assign dSP_558_b = _zz_b_4[111 : 104];
  assign dSP_559_a = loadWeight_1_weightRead_4_data[631 : 624];
  assign dSP_559_d = loadWeight_1_weightRead_4_data[759 : 752];
  assign dSP_559_b = _zz_b_4[119 : 112];
  assign dSP_560_a = loadWeight_1_weightRead_4_data[639 : 632];
  assign dSP_560_d = loadWeight_1_weightRead_4_data[767 : 760];
  assign dSP_560_b = _zz_b_4[127 : 120];
  assign dSP_561_a = loadWeight_1_weightRead_4_data[775 : 768];
  assign dSP_561_d = loadWeight_1_weightRead_4_data[903 : 896];
  assign dSP_561_b = _zz_b_4[7 : 0];
  assign dSP_562_a = loadWeight_1_weightRead_4_data[783 : 776];
  assign dSP_562_d = loadWeight_1_weightRead_4_data[911 : 904];
  assign dSP_562_b = _zz_b_4[15 : 8];
  assign dSP_563_a = loadWeight_1_weightRead_4_data[791 : 784];
  assign dSP_563_d = loadWeight_1_weightRead_4_data[919 : 912];
  assign dSP_563_b = _zz_b_4[23 : 16];
  assign dSP_564_a = loadWeight_1_weightRead_4_data[799 : 792];
  assign dSP_564_d = loadWeight_1_weightRead_4_data[927 : 920];
  assign dSP_564_b = _zz_b_4[31 : 24];
  assign dSP_565_a = loadWeight_1_weightRead_4_data[807 : 800];
  assign dSP_565_d = loadWeight_1_weightRead_4_data[935 : 928];
  assign dSP_565_b = _zz_b_4[39 : 32];
  assign dSP_566_a = loadWeight_1_weightRead_4_data[815 : 808];
  assign dSP_566_d = loadWeight_1_weightRead_4_data[943 : 936];
  assign dSP_566_b = _zz_b_4[47 : 40];
  assign dSP_567_a = loadWeight_1_weightRead_4_data[823 : 816];
  assign dSP_567_d = loadWeight_1_weightRead_4_data[951 : 944];
  assign dSP_567_b = _zz_b_4[55 : 48];
  assign dSP_568_a = loadWeight_1_weightRead_4_data[831 : 824];
  assign dSP_568_d = loadWeight_1_weightRead_4_data[959 : 952];
  assign dSP_568_b = _zz_b_4[63 : 56];
  assign dSP_569_a = loadWeight_1_weightRead_4_data[839 : 832];
  assign dSP_569_d = loadWeight_1_weightRead_4_data[967 : 960];
  assign dSP_569_b = _zz_b_4[71 : 64];
  assign dSP_570_a = loadWeight_1_weightRead_4_data[847 : 840];
  assign dSP_570_d = loadWeight_1_weightRead_4_data[975 : 968];
  assign dSP_570_b = _zz_b_4[79 : 72];
  assign dSP_571_a = loadWeight_1_weightRead_4_data[855 : 848];
  assign dSP_571_d = loadWeight_1_weightRead_4_data[983 : 976];
  assign dSP_571_b = _zz_b_4[87 : 80];
  assign dSP_572_a = loadWeight_1_weightRead_4_data[863 : 856];
  assign dSP_572_d = loadWeight_1_weightRead_4_data[991 : 984];
  assign dSP_572_b = _zz_b_4[95 : 88];
  assign dSP_573_a = loadWeight_1_weightRead_4_data[871 : 864];
  assign dSP_573_d = loadWeight_1_weightRead_4_data[999 : 992];
  assign dSP_573_b = _zz_b_4[103 : 96];
  assign dSP_574_a = loadWeight_1_weightRead_4_data[879 : 872];
  assign dSP_574_d = loadWeight_1_weightRead_4_data[1007 : 1000];
  assign dSP_574_b = _zz_b_4[111 : 104];
  assign dSP_575_a = loadWeight_1_weightRead_4_data[887 : 880];
  assign dSP_575_d = loadWeight_1_weightRead_4_data[1015 : 1008];
  assign dSP_575_b = _zz_b_4[119 : 112];
  assign dSP_576_a = loadWeight_1_weightRead_4_data[895 : 888];
  assign dSP_576_d = loadWeight_1_weightRead_4_data[1023 : 1016];
  assign dSP_576_b = _zz_b_4[127 : 120];
  assign dSP_577_a = loadWeight_1_weightRead_4_data[1031 : 1024];
  assign dSP_577_d = loadWeight_1_weightRead_4_data[1159 : 1152];
  assign dSP_577_b = _zz_b_4[7 : 0];
  assign dSP_578_a = loadWeight_1_weightRead_4_data[1039 : 1032];
  assign dSP_578_d = loadWeight_1_weightRead_4_data[1167 : 1160];
  assign dSP_578_b = _zz_b_4[15 : 8];
  assign dSP_579_a = loadWeight_1_weightRead_4_data[1047 : 1040];
  assign dSP_579_d = loadWeight_1_weightRead_4_data[1175 : 1168];
  assign dSP_579_b = _zz_b_4[23 : 16];
  assign dSP_580_a = loadWeight_1_weightRead_4_data[1055 : 1048];
  assign dSP_580_d = loadWeight_1_weightRead_4_data[1183 : 1176];
  assign dSP_580_b = _zz_b_4[31 : 24];
  assign dSP_581_a = loadWeight_1_weightRead_4_data[1063 : 1056];
  assign dSP_581_d = loadWeight_1_weightRead_4_data[1191 : 1184];
  assign dSP_581_b = _zz_b_4[39 : 32];
  assign dSP_582_a = loadWeight_1_weightRead_4_data[1071 : 1064];
  assign dSP_582_d = loadWeight_1_weightRead_4_data[1199 : 1192];
  assign dSP_582_b = _zz_b_4[47 : 40];
  assign dSP_583_a = loadWeight_1_weightRead_4_data[1079 : 1072];
  assign dSP_583_d = loadWeight_1_weightRead_4_data[1207 : 1200];
  assign dSP_583_b = _zz_b_4[55 : 48];
  assign dSP_584_a = loadWeight_1_weightRead_4_data[1087 : 1080];
  assign dSP_584_d = loadWeight_1_weightRead_4_data[1215 : 1208];
  assign dSP_584_b = _zz_b_4[63 : 56];
  assign dSP_585_a = loadWeight_1_weightRead_4_data[1095 : 1088];
  assign dSP_585_d = loadWeight_1_weightRead_4_data[1223 : 1216];
  assign dSP_585_b = _zz_b_4[71 : 64];
  assign dSP_586_a = loadWeight_1_weightRead_4_data[1103 : 1096];
  assign dSP_586_d = loadWeight_1_weightRead_4_data[1231 : 1224];
  assign dSP_586_b = _zz_b_4[79 : 72];
  assign dSP_587_a = loadWeight_1_weightRead_4_data[1111 : 1104];
  assign dSP_587_d = loadWeight_1_weightRead_4_data[1239 : 1232];
  assign dSP_587_b = _zz_b_4[87 : 80];
  assign dSP_588_a = loadWeight_1_weightRead_4_data[1119 : 1112];
  assign dSP_588_d = loadWeight_1_weightRead_4_data[1247 : 1240];
  assign dSP_588_b = _zz_b_4[95 : 88];
  assign dSP_589_a = loadWeight_1_weightRead_4_data[1127 : 1120];
  assign dSP_589_d = loadWeight_1_weightRead_4_data[1255 : 1248];
  assign dSP_589_b = _zz_b_4[103 : 96];
  assign dSP_590_a = loadWeight_1_weightRead_4_data[1135 : 1128];
  assign dSP_590_d = loadWeight_1_weightRead_4_data[1263 : 1256];
  assign dSP_590_b = _zz_b_4[111 : 104];
  assign dSP_591_a = loadWeight_1_weightRead_4_data[1143 : 1136];
  assign dSP_591_d = loadWeight_1_weightRead_4_data[1271 : 1264];
  assign dSP_591_b = _zz_b_4[119 : 112];
  assign dSP_592_a = loadWeight_1_weightRead_4_data[1151 : 1144];
  assign dSP_592_d = loadWeight_1_weightRead_4_data[1279 : 1272];
  assign dSP_592_b = _zz_b_4[127 : 120];
  assign dSP_593_a = loadWeight_1_weightRead_4_data[1287 : 1280];
  assign dSP_593_d = loadWeight_1_weightRead_4_data[1415 : 1408];
  assign dSP_593_b = _zz_b_4[7 : 0];
  assign dSP_594_a = loadWeight_1_weightRead_4_data[1295 : 1288];
  assign dSP_594_d = loadWeight_1_weightRead_4_data[1423 : 1416];
  assign dSP_594_b = _zz_b_4[15 : 8];
  assign dSP_595_a = loadWeight_1_weightRead_4_data[1303 : 1296];
  assign dSP_595_d = loadWeight_1_weightRead_4_data[1431 : 1424];
  assign dSP_595_b = _zz_b_4[23 : 16];
  assign dSP_596_a = loadWeight_1_weightRead_4_data[1311 : 1304];
  assign dSP_596_d = loadWeight_1_weightRead_4_data[1439 : 1432];
  assign dSP_596_b = _zz_b_4[31 : 24];
  assign dSP_597_a = loadWeight_1_weightRead_4_data[1319 : 1312];
  assign dSP_597_d = loadWeight_1_weightRead_4_data[1447 : 1440];
  assign dSP_597_b = _zz_b_4[39 : 32];
  assign dSP_598_a = loadWeight_1_weightRead_4_data[1327 : 1320];
  assign dSP_598_d = loadWeight_1_weightRead_4_data[1455 : 1448];
  assign dSP_598_b = _zz_b_4[47 : 40];
  assign dSP_599_a = loadWeight_1_weightRead_4_data[1335 : 1328];
  assign dSP_599_d = loadWeight_1_weightRead_4_data[1463 : 1456];
  assign dSP_599_b = _zz_b_4[55 : 48];
  assign dSP_600_a = loadWeight_1_weightRead_4_data[1343 : 1336];
  assign dSP_600_d = loadWeight_1_weightRead_4_data[1471 : 1464];
  assign dSP_600_b = _zz_b_4[63 : 56];
  assign dSP_601_a = loadWeight_1_weightRead_4_data[1351 : 1344];
  assign dSP_601_d = loadWeight_1_weightRead_4_data[1479 : 1472];
  assign dSP_601_b = _zz_b_4[71 : 64];
  assign dSP_602_a = loadWeight_1_weightRead_4_data[1359 : 1352];
  assign dSP_602_d = loadWeight_1_weightRead_4_data[1487 : 1480];
  assign dSP_602_b = _zz_b_4[79 : 72];
  assign dSP_603_a = loadWeight_1_weightRead_4_data[1367 : 1360];
  assign dSP_603_d = loadWeight_1_weightRead_4_data[1495 : 1488];
  assign dSP_603_b = _zz_b_4[87 : 80];
  assign dSP_604_a = loadWeight_1_weightRead_4_data[1375 : 1368];
  assign dSP_604_d = loadWeight_1_weightRead_4_data[1503 : 1496];
  assign dSP_604_b = _zz_b_4[95 : 88];
  assign dSP_605_a = loadWeight_1_weightRead_4_data[1383 : 1376];
  assign dSP_605_d = loadWeight_1_weightRead_4_data[1511 : 1504];
  assign dSP_605_b = _zz_b_4[103 : 96];
  assign dSP_606_a = loadWeight_1_weightRead_4_data[1391 : 1384];
  assign dSP_606_d = loadWeight_1_weightRead_4_data[1519 : 1512];
  assign dSP_606_b = _zz_b_4[111 : 104];
  assign dSP_607_a = loadWeight_1_weightRead_4_data[1399 : 1392];
  assign dSP_607_d = loadWeight_1_weightRead_4_data[1527 : 1520];
  assign dSP_607_b = _zz_b_4[119 : 112];
  assign dSP_608_a = loadWeight_1_weightRead_4_data[1407 : 1400];
  assign dSP_608_d = loadWeight_1_weightRead_4_data[1535 : 1528];
  assign dSP_608_b = _zz_b_4[127 : 120];
  assign dSP_609_a = loadWeight_1_weightRead_4_data[1543 : 1536];
  assign dSP_609_d = loadWeight_1_weightRead_4_data[1671 : 1664];
  assign dSP_609_b = _zz_b_4[7 : 0];
  assign dSP_610_a = loadWeight_1_weightRead_4_data[1551 : 1544];
  assign dSP_610_d = loadWeight_1_weightRead_4_data[1679 : 1672];
  assign dSP_610_b = _zz_b_4[15 : 8];
  assign dSP_611_a = loadWeight_1_weightRead_4_data[1559 : 1552];
  assign dSP_611_d = loadWeight_1_weightRead_4_data[1687 : 1680];
  assign dSP_611_b = _zz_b_4[23 : 16];
  assign dSP_612_a = loadWeight_1_weightRead_4_data[1567 : 1560];
  assign dSP_612_d = loadWeight_1_weightRead_4_data[1695 : 1688];
  assign dSP_612_b = _zz_b_4[31 : 24];
  assign dSP_613_a = loadWeight_1_weightRead_4_data[1575 : 1568];
  assign dSP_613_d = loadWeight_1_weightRead_4_data[1703 : 1696];
  assign dSP_613_b = _zz_b_4[39 : 32];
  assign dSP_614_a = loadWeight_1_weightRead_4_data[1583 : 1576];
  assign dSP_614_d = loadWeight_1_weightRead_4_data[1711 : 1704];
  assign dSP_614_b = _zz_b_4[47 : 40];
  assign dSP_615_a = loadWeight_1_weightRead_4_data[1591 : 1584];
  assign dSP_615_d = loadWeight_1_weightRead_4_data[1719 : 1712];
  assign dSP_615_b = _zz_b_4[55 : 48];
  assign dSP_616_a = loadWeight_1_weightRead_4_data[1599 : 1592];
  assign dSP_616_d = loadWeight_1_weightRead_4_data[1727 : 1720];
  assign dSP_616_b = _zz_b_4[63 : 56];
  assign dSP_617_a = loadWeight_1_weightRead_4_data[1607 : 1600];
  assign dSP_617_d = loadWeight_1_weightRead_4_data[1735 : 1728];
  assign dSP_617_b = _zz_b_4[71 : 64];
  assign dSP_618_a = loadWeight_1_weightRead_4_data[1615 : 1608];
  assign dSP_618_d = loadWeight_1_weightRead_4_data[1743 : 1736];
  assign dSP_618_b = _zz_b_4[79 : 72];
  assign dSP_619_a = loadWeight_1_weightRead_4_data[1623 : 1616];
  assign dSP_619_d = loadWeight_1_weightRead_4_data[1751 : 1744];
  assign dSP_619_b = _zz_b_4[87 : 80];
  assign dSP_620_a = loadWeight_1_weightRead_4_data[1631 : 1624];
  assign dSP_620_d = loadWeight_1_weightRead_4_data[1759 : 1752];
  assign dSP_620_b = _zz_b_4[95 : 88];
  assign dSP_621_a = loadWeight_1_weightRead_4_data[1639 : 1632];
  assign dSP_621_d = loadWeight_1_weightRead_4_data[1767 : 1760];
  assign dSP_621_b = _zz_b_4[103 : 96];
  assign dSP_622_a = loadWeight_1_weightRead_4_data[1647 : 1640];
  assign dSP_622_d = loadWeight_1_weightRead_4_data[1775 : 1768];
  assign dSP_622_b = _zz_b_4[111 : 104];
  assign dSP_623_a = loadWeight_1_weightRead_4_data[1655 : 1648];
  assign dSP_623_d = loadWeight_1_weightRead_4_data[1783 : 1776];
  assign dSP_623_b = _zz_b_4[119 : 112];
  assign dSP_624_a = loadWeight_1_weightRead_4_data[1663 : 1656];
  assign dSP_624_d = loadWeight_1_weightRead_4_data[1791 : 1784];
  assign dSP_624_b = _zz_b_4[127 : 120];
  assign dSP_625_a = loadWeight_1_weightRead_4_data[1799 : 1792];
  assign dSP_625_d = loadWeight_1_weightRead_4_data[1927 : 1920];
  assign dSP_625_b = _zz_b_4[7 : 0];
  assign dSP_626_a = loadWeight_1_weightRead_4_data[1807 : 1800];
  assign dSP_626_d = loadWeight_1_weightRead_4_data[1935 : 1928];
  assign dSP_626_b = _zz_b_4[15 : 8];
  assign dSP_627_a = loadWeight_1_weightRead_4_data[1815 : 1808];
  assign dSP_627_d = loadWeight_1_weightRead_4_data[1943 : 1936];
  assign dSP_627_b = _zz_b_4[23 : 16];
  assign dSP_628_a = loadWeight_1_weightRead_4_data[1823 : 1816];
  assign dSP_628_d = loadWeight_1_weightRead_4_data[1951 : 1944];
  assign dSP_628_b = _zz_b_4[31 : 24];
  assign dSP_629_a = loadWeight_1_weightRead_4_data[1831 : 1824];
  assign dSP_629_d = loadWeight_1_weightRead_4_data[1959 : 1952];
  assign dSP_629_b = _zz_b_4[39 : 32];
  assign dSP_630_a = loadWeight_1_weightRead_4_data[1839 : 1832];
  assign dSP_630_d = loadWeight_1_weightRead_4_data[1967 : 1960];
  assign dSP_630_b = _zz_b_4[47 : 40];
  assign dSP_631_a = loadWeight_1_weightRead_4_data[1847 : 1840];
  assign dSP_631_d = loadWeight_1_weightRead_4_data[1975 : 1968];
  assign dSP_631_b = _zz_b_4[55 : 48];
  assign dSP_632_a = loadWeight_1_weightRead_4_data[1855 : 1848];
  assign dSP_632_d = loadWeight_1_weightRead_4_data[1983 : 1976];
  assign dSP_632_b = _zz_b_4[63 : 56];
  assign dSP_633_a = loadWeight_1_weightRead_4_data[1863 : 1856];
  assign dSP_633_d = loadWeight_1_weightRead_4_data[1991 : 1984];
  assign dSP_633_b = _zz_b_4[71 : 64];
  assign dSP_634_a = loadWeight_1_weightRead_4_data[1871 : 1864];
  assign dSP_634_d = loadWeight_1_weightRead_4_data[1999 : 1992];
  assign dSP_634_b = _zz_b_4[79 : 72];
  assign dSP_635_a = loadWeight_1_weightRead_4_data[1879 : 1872];
  assign dSP_635_d = loadWeight_1_weightRead_4_data[2007 : 2000];
  assign dSP_635_b = _zz_b_4[87 : 80];
  assign dSP_636_a = loadWeight_1_weightRead_4_data[1887 : 1880];
  assign dSP_636_d = loadWeight_1_weightRead_4_data[2015 : 2008];
  assign dSP_636_b = _zz_b_4[95 : 88];
  assign dSP_637_a = loadWeight_1_weightRead_4_data[1895 : 1888];
  assign dSP_637_d = loadWeight_1_weightRead_4_data[2023 : 2016];
  assign dSP_637_b = _zz_b_4[103 : 96];
  assign dSP_638_a = loadWeight_1_weightRead_4_data[1903 : 1896];
  assign dSP_638_d = loadWeight_1_weightRead_4_data[2031 : 2024];
  assign dSP_638_b = _zz_b_4[111 : 104];
  assign dSP_639_a = loadWeight_1_weightRead_4_data[1911 : 1904];
  assign dSP_639_d = loadWeight_1_weightRead_4_data[2039 : 2032];
  assign dSP_639_b = _zz_b_4[119 : 112];
  assign dSP_640_a = loadWeight_1_weightRead_4_data[1919 : 1912];
  assign dSP_640_d = loadWeight_1_weightRead_4_data[2047 : 2040];
  assign dSP_640_b = _zz_b_4[127 : 120];
  assign dSP_641_a = loadWeight_1_weightRead_5_data[7 : 0];
  assign dSP_641_d = loadWeight_1_weightRead_5_data[135 : 128];
  assign dSP_641_b = _zz_b_5[7 : 0];
  assign dSP_642_a = loadWeight_1_weightRead_5_data[15 : 8];
  assign dSP_642_d = loadWeight_1_weightRead_5_data[143 : 136];
  assign dSP_642_b = _zz_b_5[15 : 8];
  assign dSP_643_a = loadWeight_1_weightRead_5_data[23 : 16];
  assign dSP_643_d = loadWeight_1_weightRead_5_data[151 : 144];
  assign dSP_643_b = _zz_b_5[23 : 16];
  assign dSP_644_a = loadWeight_1_weightRead_5_data[31 : 24];
  assign dSP_644_d = loadWeight_1_weightRead_5_data[159 : 152];
  assign dSP_644_b = _zz_b_5[31 : 24];
  assign dSP_645_a = loadWeight_1_weightRead_5_data[39 : 32];
  assign dSP_645_d = loadWeight_1_weightRead_5_data[167 : 160];
  assign dSP_645_b = _zz_b_5[39 : 32];
  assign dSP_646_a = loadWeight_1_weightRead_5_data[47 : 40];
  assign dSP_646_d = loadWeight_1_weightRead_5_data[175 : 168];
  assign dSP_646_b = _zz_b_5[47 : 40];
  assign dSP_647_a = loadWeight_1_weightRead_5_data[55 : 48];
  assign dSP_647_d = loadWeight_1_weightRead_5_data[183 : 176];
  assign dSP_647_b = _zz_b_5[55 : 48];
  assign dSP_648_a = loadWeight_1_weightRead_5_data[63 : 56];
  assign dSP_648_d = loadWeight_1_weightRead_5_data[191 : 184];
  assign dSP_648_b = _zz_b_5[63 : 56];
  assign dSP_649_a = loadWeight_1_weightRead_5_data[71 : 64];
  assign dSP_649_d = loadWeight_1_weightRead_5_data[199 : 192];
  assign dSP_649_b = _zz_b_5[71 : 64];
  assign dSP_650_a = loadWeight_1_weightRead_5_data[79 : 72];
  assign dSP_650_d = loadWeight_1_weightRead_5_data[207 : 200];
  assign dSP_650_b = _zz_b_5[79 : 72];
  assign dSP_651_a = loadWeight_1_weightRead_5_data[87 : 80];
  assign dSP_651_d = loadWeight_1_weightRead_5_data[215 : 208];
  assign dSP_651_b = _zz_b_5[87 : 80];
  assign dSP_652_a = loadWeight_1_weightRead_5_data[95 : 88];
  assign dSP_652_d = loadWeight_1_weightRead_5_data[223 : 216];
  assign dSP_652_b = _zz_b_5[95 : 88];
  assign dSP_653_a = loadWeight_1_weightRead_5_data[103 : 96];
  assign dSP_653_d = loadWeight_1_weightRead_5_data[231 : 224];
  assign dSP_653_b = _zz_b_5[103 : 96];
  assign dSP_654_a = loadWeight_1_weightRead_5_data[111 : 104];
  assign dSP_654_d = loadWeight_1_weightRead_5_data[239 : 232];
  assign dSP_654_b = _zz_b_5[111 : 104];
  assign dSP_655_a = loadWeight_1_weightRead_5_data[119 : 112];
  assign dSP_655_d = loadWeight_1_weightRead_5_data[247 : 240];
  assign dSP_655_b = _zz_b_5[119 : 112];
  assign dSP_656_a = loadWeight_1_weightRead_5_data[127 : 120];
  assign dSP_656_d = loadWeight_1_weightRead_5_data[255 : 248];
  assign dSP_656_b = _zz_b_5[127 : 120];
  assign dSP_657_a = loadWeight_1_weightRead_5_data[263 : 256];
  assign dSP_657_d = loadWeight_1_weightRead_5_data[391 : 384];
  assign dSP_657_b = _zz_b_5[7 : 0];
  assign dSP_658_a = loadWeight_1_weightRead_5_data[271 : 264];
  assign dSP_658_d = loadWeight_1_weightRead_5_data[399 : 392];
  assign dSP_658_b = _zz_b_5[15 : 8];
  assign dSP_659_a = loadWeight_1_weightRead_5_data[279 : 272];
  assign dSP_659_d = loadWeight_1_weightRead_5_data[407 : 400];
  assign dSP_659_b = _zz_b_5[23 : 16];
  assign dSP_660_a = loadWeight_1_weightRead_5_data[287 : 280];
  assign dSP_660_d = loadWeight_1_weightRead_5_data[415 : 408];
  assign dSP_660_b = _zz_b_5[31 : 24];
  assign dSP_661_a = loadWeight_1_weightRead_5_data[295 : 288];
  assign dSP_661_d = loadWeight_1_weightRead_5_data[423 : 416];
  assign dSP_661_b = _zz_b_5[39 : 32];
  assign dSP_662_a = loadWeight_1_weightRead_5_data[303 : 296];
  assign dSP_662_d = loadWeight_1_weightRead_5_data[431 : 424];
  assign dSP_662_b = _zz_b_5[47 : 40];
  assign dSP_663_a = loadWeight_1_weightRead_5_data[311 : 304];
  assign dSP_663_d = loadWeight_1_weightRead_5_data[439 : 432];
  assign dSP_663_b = _zz_b_5[55 : 48];
  assign dSP_664_a = loadWeight_1_weightRead_5_data[319 : 312];
  assign dSP_664_d = loadWeight_1_weightRead_5_data[447 : 440];
  assign dSP_664_b = _zz_b_5[63 : 56];
  assign dSP_665_a = loadWeight_1_weightRead_5_data[327 : 320];
  assign dSP_665_d = loadWeight_1_weightRead_5_data[455 : 448];
  assign dSP_665_b = _zz_b_5[71 : 64];
  assign dSP_666_a = loadWeight_1_weightRead_5_data[335 : 328];
  assign dSP_666_d = loadWeight_1_weightRead_5_data[463 : 456];
  assign dSP_666_b = _zz_b_5[79 : 72];
  assign dSP_667_a = loadWeight_1_weightRead_5_data[343 : 336];
  assign dSP_667_d = loadWeight_1_weightRead_5_data[471 : 464];
  assign dSP_667_b = _zz_b_5[87 : 80];
  assign dSP_668_a = loadWeight_1_weightRead_5_data[351 : 344];
  assign dSP_668_d = loadWeight_1_weightRead_5_data[479 : 472];
  assign dSP_668_b = _zz_b_5[95 : 88];
  assign dSP_669_a = loadWeight_1_weightRead_5_data[359 : 352];
  assign dSP_669_d = loadWeight_1_weightRead_5_data[487 : 480];
  assign dSP_669_b = _zz_b_5[103 : 96];
  assign dSP_670_a = loadWeight_1_weightRead_5_data[367 : 360];
  assign dSP_670_d = loadWeight_1_weightRead_5_data[495 : 488];
  assign dSP_670_b = _zz_b_5[111 : 104];
  assign dSP_671_a = loadWeight_1_weightRead_5_data[375 : 368];
  assign dSP_671_d = loadWeight_1_weightRead_5_data[503 : 496];
  assign dSP_671_b = _zz_b_5[119 : 112];
  assign dSP_672_a = loadWeight_1_weightRead_5_data[383 : 376];
  assign dSP_672_d = loadWeight_1_weightRead_5_data[511 : 504];
  assign dSP_672_b = _zz_b_5[127 : 120];
  assign dSP_673_a = loadWeight_1_weightRead_5_data[519 : 512];
  assign dSP_673_d = loadWeight_1_weightRead_5_data[647 : 640];
  assign dSP_673_b = _zz_b_5[7 : 0];
  assign dSP_674_a = loadWeight_1_weightRead_5_data[527 : 520];
  assign dSP_674_d = loadWeight_1_weightRead_5_data[655 : 648];
  assign dSP_674_b = _zz_b_5[15 : 8];
  assign dSP_675_a = loadWeight_1_weightRead_5_data[535 : 528];
  assign dSP_675_d = loadWeight_1_weightRead_5_data[663 : 656];
  assign dSP_675_b = _zz_b_5[23 : 16];
  assign dSP_676_a = loadWeight_1_weightRead_5_data[543 : 536];
  assign dSP_676_d = loadWeight_1_weightRead_5_data[671 : 664];
  assign dSP_676_b = _zz_b_5[31 : 24];
  assign dSP_677_a = loadWeight_1_weightRead_5_data[551 : 544];
  assign dSP_677_d = loadWeight_1_weightRead_5_data[679 : 672];
  assign dSP_677_b = _zz_b_5[39 : 32];
  assign dSP_678_a = loadWeight_1_weightRead_5_data[559 : 552];
  assign dSP_678_d = loadWeight_1_weightRead_5_data[687 : 680];
  assign dSP_678_b = _zz_b_5[47 : 40];
  assign dSP_679_a = loadWeight_1_weightRead_5_data[567 : 560];
  assign dSP_679_d = loadWeight_1_weightRead_5_data[695 : 688];
  assign dSP_679_b = _zz_b_5[55 : 48];
  assign dSP_680_a = loadWeight_1_weightRead_5_data[575 : 568];
  assign dSP_680_d = loadWeight_1_weightRead_5_data[703 : 696];
  assign dSP_680_b = _zz_b_5[63 : 56];
  assign dSP_681_a = loadWeight_1_weightRead_5_data[583 : 576];
  assign dSP_681_d = loadWeight_1_weightRead_5_data[711 : 704];
  assign dSP_681_b = _zz_b_5[71 : 64];
  assign dSP_682_a = loadWeight_1_weightRead_5_data[591 : 584];
  assign dSP_682_d = loadWeight_1_weightRead_5_data[719 : 712];
  assign dSP_682_b = _zz_b_5[79 : 72];
  assign dSP_683_a = loadWeight_1_weightRead_5_data[599 : 592];
  assign dSP_683_d = loadWeight_1_weightRead_5_data[727 : 720];
  assign dSP_683_b = _zz_b_5[87 : 80];
  assign dSP_684_a = loadWeight_1_weightRead_5_data[607 : 600];
  assign dSP_684_d = loadWeight_1_weightRead_5_data[735 : 728];
  assign dSP_684_b = _zz_b_5[95 : 88];
  assign dSP_685_a = loadWeight_1_weightRead_5_data[615 : 608];
  assign dSP_685_d = loadWeight_1_weightRead_5_data[743 : 736];
  assign dSP_685_b = _zz_b_5[103 : 96];
  assign dSP_686_a = loadWeight_1_weightRead_5_data[623 : 616];
  assign dSP_686_d = loadWeight_1_weightRead_5_data[751 : 744];
  assign dSP_686_b = _zz_b_5[111 : 104];
  assign dSP_687_a = loadWeight_1_weightRead_5_data[631 : 624];
  assign dSP_687_d = loadWeight_1_weightRead_5_data[759 : 752];
  assign dSP_687_b = _zz_b_5[119 : 112];
  assign dSP_688_a = loadWeight_1_weightRead_5_data[639 : 632];
  assign dSP_688_d = loadWeight_1_weightRead_5_data[767 : 760];
  assign dSP_688_b = _zz_b_5[127 : 120];
  assign dSP_689_a = loadWeight_1_weightRead_5_data[775 : 768];
  assign dSP_689_d = loadWeight_1_weightRead_5_data[903 : 896];
  assign dSP_689_b = _zz_b_5[7 : 0];
  assign dSP_690_a = loadWeight_1_weightRead_5_data[783 : 776];
  assign dSP_690_d = loadWeight_1_weightRead_5_data[911 : 904];
  assign dSP_690_b = _zz_b_5[15 : 8];
  assign dSP_691_a = loadWeight_1_weightRead_5_data[791 : 784];
  assign dSP_691_d = loadWeight_1_weightRead_5_data[919 : 912];
  assign dSP_691_b = _zz_b_5[23 : 16];
  assign dSP_692_a = loadWeight_1_weightRead_5_data[799 : 792];
  assign dSP_692_d = loadWeight_1_weightRead_5_data[927 : 920];
  assign dSP_692_b = _zz_b_5[31 : 24];
  assign dSP_693_a = loadWeight_1_weightRead_5_data[807 : 800];
  assign dSP_693_d = loadWeight_1_weightRead_5_data[935 : 928];
  assign dSP_693_b = _zz_b_5[39 : 32];
  assign dSP_694_a = loadWeight_1_weightRead_5_data[815 : 808];
  assign dSP_694_d = loadWeight_1_weightRead_5_data[943 : 936];
  assign dSP_694_b = _zz_b_5[47 : 40];
  assign dSP_695_a = loadWeight_1_weightRead_5_data[823 : 816];
  assign dSP_695_d = loadWeight_1_weightRead_5_data[951 : 944];
  assign dSP_695_b = _zz_b_5[55 : 48];
  assign dSP_696_a = loadWeight_1_weightRead_5_data[831 : 824];
  assign dSP_696_d = loadWeight_1_weightRead_5_data[959 : 952];
  assign dSP_696_b = _zz_b_5[63 : 56];
  assign dSP_697_a = loadWeight_1_weightRead_5_data[839 : 832];
  assign dSP_697_d = loadWeight_1_weightRead_5_data[967 : 960];
  assign dSP_697_b = _zz_b_5[71 : 64];
  assign dSP_698_a = loadWeight_1_weightRead_5_data[847 : 840];
  assign dSP_698_d = loadWeight_1_weightRead_5_data[975 : 968];
  assign dSP_698_b = _zz_b_5[79 : 72];
  assign dSP_699_a = loadWeight_1_weightRead_5_data[855 : 848];
  assign dSP_699_d = loadWeight_1_weightRead_5_data[983 : 976];
  assign dSP_699_b = _zz_b_5[87 : 80];
  assign dSP_700_a = loadWeight_1_weightRead_5_data[863 : 856];
  assign dSP_700_d = loadWeight_1_weightRead_5_data[991 : 984];
  assign dSP_700_b = _zz_b_5[95 : 88];
  assign dSP_701_a = loadWeight_1_weightRead_5_data[871 : 864];
  assign dSP_701_d = loadWeight_1_weightRead_5_data[999 : 992];
  assign dSP_701_b = _zz_b_5[103 : 96];
  assign dSP_702_a = loadWeight_1_weightRead_5_data[879 : 872];
  assign dSP_702_d = loadWeight_1_weightRead_5_data[1007 : 1000];
  assign dSP_702_b = _zz_b_5[111 : 104];
  assign dSP_703_a = loadWeight_1_weightRead_5_data[887 : 880];
  assign dSP_703_d = loadWeight_1_weightRead_5_data[1015 : 1008];
  assign dSP_703_b = _zz_b_5[119 : 112];
  assign dSP_704_a = loadWeight_1_weightRead_5_data[895 : 888];
  assign dSP_704_d = loadWeight_1_weightRead_5_data[1023 : 1016];
  assign dSP_704_b = _zz_b_5[127 : 120];
  assign dSP_705_a = loadWeight_1_weightRead_5_data[1031 : 1024];
  assign dSP_705_d = loadWeight_1_weightRead_5_data[1159 : 1152];
  assign dSP_705_b = _zz_b_5[7 : 0];
  assign dSP_706_a = loadWeight_1_weightRead_5_data[1039 : 1032];
  assign dSP_706_d = loadWeight_1_weightRead_5_data[1167 : 1160];
  assign dSP_706_b = _zz_b_5[15 : 8];
  assign dSP_707_a = loadWeight_1_weightRead_5_data[1047 : 1040];
  assign dSP_707_d = loadWeight_1_weightRead_5_data[1175 : 1168];
  assign dSP_707_b = _zz_b_5[23 : 16];
  assign dSP_708_a = loadWeight_1_weightRead_5_data[1055 : 1048];
  assign dSP_708_d = loadWeight_1_weightRead_5_data[1183 : 1176];
  assign dSP_708_b = _zz_b_5[31 : 24];
  assign dSP_709_a = loadWeight_1_weightRead_5_data[1063 : 1056];
  assign dSP_709_d = loadWeight_1_weightRead_5_data[1191 : 1184];
  assign dSP_709_b = _zz_b_5[39 : 32];
  assign dSP_710_a = loadWeight_1_weightRead_5_data[1071 : 1064];
  assign dSP_710_d = loadWeight_1_weightRead_5_data[1199 : 1192];
  assign dSP_710_b = _zz_b_5[47 : 40];
  assign dSP_711_a = loadWeight_1_weightRead_5_data[1079 : 1072];
  assign dSP_711_d = loadWeight_1_weightRead_5_data[1207 : 1200];
  assign dSP_711_b = _zz_b_5[55 : 48];
  assign dSP_712_a = loadWeight_1_weightRead_5_data[1087 : 1080];
  assign dSP_712_d = loadWeight_1_weightRead_5_data[1215 : 1208];
  assign dSP_712_b = _zz_b_5[63 : 56];
  assign dSP_713_a = loadWeight_1_weightRead_5_data[1095 : 1088];
  assign dSP_713_d = loadWeight_1_weightRead_5_data[1223 : 1216];
  assign dSP_713_b = _zz_b_5[71 : 64];
  assign dSP_714_a = loadWeight_1_weightRead_5_data[1103 : 1096];
  assign dSP_714_d = loadWeight_1_weightRead_5_data[1231 : 1224];
  assign dSP_714_b = _zz_b_5[79 : 72];
  assign dSP_715_a = loadWeight_1_weightRead_5_data[1111 : 1104];
  assign dSP_715_d = loadWeight_1_weightRead_5_data[1239 : 1232];
  assign dSP_715_b = _zz_b_5[87 : 80];
  assign dSP_716_a = loadWeight_1_weightRead_5_data[1119 : 1112];
  assign dSP_716_d = loadWeight_1_weightRead_5_data[1247 : 1240];
  assign dSP_716_b = _zz_b_5[95 : 88];
  assign dSP_717_a = loadWeight_1_weightRead_5_data[1127 : 1120];
  assign dSP_717_d = loadWeight_1_weightRead_5_data[1255 : 1248];
  assign dSP_717_b = _zz_b_5[103 : 96];
  assign dSP_718_a = loadWeight_1_weightRead_5_data[1135 : 1128];
  assign dSP_718_d = loadWeight_1_weightRead_5_data[1263 : 1256];
  assign dSP_718_b = _zz_b_5[111 : 104];
  assign dSP_719_a = loadWeight_1_weightRead_5_data[1143 : 1136];
  assign dSP_719_d = loadWeight_1_weightRead_5_data[1271 : 1264];
  assign dSP_719_b = _zz_b_5[119 : 112];
  assign dSP_720_a = loadWeight_1_weightRead_5_data[1151 : 1144];
  assign dSP_720_d = loadWeight_1_weightRead_5_data[1279 : 1272];
  assign dSP_720_b = _zz_b_5[127 : 120];
  assign dSP_721_a = loadWeight_1_weightRead_5_data[1287 : 1280];
  assign dSP_721_d = loadWeight_1_weightRead_5_data[1415 : 1408];
  assign dSP_721_b = _zz_b_5[7 : 0];
  assign dSP_722_a = loadWeight_1_weightRead_5_data[1295 : 1288];
  assign dSP_722_d = loadWeight_1_weightRead_5_data[1423 : 1416];
  assign dSP_722_b = _zz_b_5[15 : 8];
  assign dSP_723_a = loadWeight_1_weightRead_5_data[1303 : 1296];
  assign dSP_723_d = loadWeight_1_weightRead_5_data[1431 : 1424];
  assign dSP_723_b = _zz_b_5[23 : 16];
  assign dSP_724_a = loadWeight_1_weightRead_5_data[1311 : 1304];
  assign dSP_724_d = loadWeight_1_weightRead_5_data[1439 : 1432];
  assign dSP_724_b = _zz_b_5[31 : 24];
  assign dSP_725_a = loadWeight_1_weightRead_5_data[1319 : 1312];
  assign dSP_725_d = loadWeight_1_weightRead_5_data[1447 : 1440];
  assign dSP_725_b = _zz_b_5[39 : 32];
  assign dSP_726_a = loadWeight_1_weightRead_5_data[1327 : 1320];
  assign dSP_726_d = loadWeight_1_weightRead_5_data[1455 : 1448];
  assign dSP_726_b = _zz_b_5[47 : 40];
  assign dSP_727_a = loadWeight_1_weightRead_5_data[1335 : 1328];
  assign dSP_727_d = loadWeight_1_weightRead_5_data[1463 : 1456];
  assign dSP_727_b = _zz_b_5[55 : 48];
  assign dSP_728_a = loadWeight_1_weightRead_5_data[1343 : 1336];
  assign dSP_728_d = loadWeight_1_weightRead_5_data[1471 : 1464];
  assign dSP_728_b = _zz_b_5[63 : 56];
  assign dSP_729_a = loadWeight_1_weightRead_5_data[1351 : 1344];
  assign dSP_729_d = loadWeight_1_weightRead_5_data[1479 : 1472];
  assign dSP_729_b = _zz_b_5[71 : 64];
  assign dSP_730_a = loadWeight_1_weightRead_5_data[1359 : 1352];
  assign dSP_730_d = loadWeight_1_weightRead_5_data[1487 : 1480];
  assign dSP_730_b = _zz_b_5[79 : 72];
  assign dSP_731_a = loadWeight_1_weightRead_5_data[1367 : 1360];
  assign dSP_731_d = loadWeight_1_weightRead_5_data[1495 : 1488];
  assign dSP_731_b = _zz_b_5[87 : 80];
  assign dSP_732_a = loadWeight_1_weightRead_5_data[1375 : 1368];
  assign dSP_732_d = loadWeight_1_weightRead_5_data[1503 : 1496];
  assign dSP_732_b = _zz_b_5[95 : 88];
  assign dSP_733_a = loadWeight_1_weightRead_5_data[1383 : 1376];
  assign dSP_733_d = loadWeight_1_weightRead_5_data[1511 : 1504];
  assign dSP_733_b = _zz_b_5[103 : 96];
  assign dSP_734_a = loadWeight_1_weightRead_5_data[1391 : 1384];
  assign dSP_734_d = loadWeight_1_weightRead_5_data[1519 : 1512];
  assign dSP_734_b = _zz_b_5[111 : 104];
  assign dSP_735_a = loadWeight_1_weightRead_5_data[1399 : 1392];
  assign dSP_735_d = loadWeight_1_weightRead_5_data[1527 : 1520];
  assign dSP_735_b = _zz_b_5[119 : 112];
  assign dSP_736_a = loadWeight_1_weightRead_5_data[1407 : 1400];
  assign dSP_736_d = loadWeight_1_weightRead_5_data[1535 : 1528];
  assign dSP_736_b = _zz_b_5[127 : 120];
  assign dSP_737_a = loadWeight_1_weightRead_5_data[1543 : 1536];
  assign dSP_737_d = loadWeight_1_weightRead_5_data[1671 : 1664];
  assign dSP_737_b = _zz_b_5[7 : 0];
  assign dSP_738_a = loadWeight_1_weightRead_5_data[1551 : 1544];
  assign dSP_738_d = loadWeight_1_weightRead_5_data[1679 : 1672];
  assign dSP_738_b = _zz_b_5[15 : 8];
  assign dSP_739_a = loadWeight_1_weightRead_5_data[1559 : 1552];
  assign dSP_739_d = loadWeight_1_weightRead_5_data[1687 : 1680];
  assign dSP_739_b = _zz_b_5[23 : 16];
  assign dSP_740_a = loadWeight_1_weightRead_5_data[1567 : 1560];
  assign dSP_740_d = loadWeight_1_weightRead_5_data[1695 : 1688];
  assign dSP_740_b = _zz_b_5[31 : 24];
  assign dSP_741_a = loadWeight_1_weightRead_5_data[1575 : 1568];
  assign dSP_741_d = loadWeight_1_weightRead_5_data[1703 : 1696];
  assign dSP_741_b = _zz_b_5[39 : 32];
  assign dSP_742_a = loadWeight_1_weightRead_5_data[1583 : 1576];
  assign dSP_742_d = loadWeight_1_weightRead_5_data[1711 : 1704];
  assign dSP_742_b = _zz_b_5[47 : 40];
  assign dSP_743_a = loadWeight_1_weightRead_5_data[1591 : 1584];
  assign dSP_743_d = loadWeight_1_weightRead_5_data[1719 : 1712];
  assign dSP_743_b = _zz_b_5[55 : 48];
  assign dSP_744_a = loadWeight_1_weightRead_5_data[1599 : 1592];
  assign dSP_744_d = loadWeight_1_weightRead_5_data[1727 : 1720];
  assign dSP_744_b = _zz_b_5[63 : 56];
  assign dSP_745_a = loadWeight_1_weightRead_5_data[1607 : 1600];
  assign dSP_745_d = loadWeight_1_weightRead_5_data[1735 : 1728];
  assign dSP_745_b = _zz_b_5[71 : 64];
  assign dSP_746_a = loadWeight_1_weightRead_5_data[1615 : 1608];
  assign dSP_746_d = loadWeight_1_weightRead_5_data[1743 : 1736];
  assign dSP_746_b = _zz_b_5[79 : 72];
  assign dSP_747_a = loadWeight_1_weightRead_5_data[1623 : 1616];
  assign dSP_747_d = loadWeight_1_weightRead_5_data[1751 : 1744];
  assign dSP_747_b = _zz_b_5[87 : 80];
  assign dSP_748_a = loadWeight_1_weightRead_5_data[1631 : 1624];
  assign dSP_748_d = loadWeight_1_weightRead_5_data[1759 : 1752];
  assign dSP_748_b = _zz_b_5[95 : 88];
  assign dSP_749_a = loadWeight_1_weightRead_5_data[1639 : 1632];
  assign dSP_749_d = loadWeight_1_weightRead_5_data[1767 : 1760];
  assign dSP_749_b = _zz_b_5[103 : 96];
  assign dSP_750_a = loadWeight_1_weightRead_5_data[1647 : 1640];
  assign dSP_750_d = loadWeight_1_weightRead_5_data[1775 : 1768];
  assign dSP_750_b = _zz_b_5[111 : 104];
  assign dSP_751_a = loadWeight_1_weightRead_5_data[1655 : 1648];
  assign dSP_751_d = loadWeight_1_weightRead_5_data[1783 : 1776];
  assign dSP_751_b = _zz_b_5[119 : 112];
  assign dSP_752_a = loadWeight_1_weightRead_5_data[1663 : 1656];
  assign dSP_752_d = loadWeight_1_weightRead_5_data[1791 : 1784];
  assign dSP_752_b = _zz_b_5[127 : 120];
  assign dSP_753_a = loadWeight_1_weightRead_5_data[1799 : 1792];
  assign dSP_753_d = loadWeight_1_weightRead_5_data[1927 : 1920];
  assign dSP_753_b = _zz_b_5[7 : 0];
  assign dSP_754_a = loadWeight_1_weightRead_5_data[1807 : 1800];
  assign dSP_754_d = loadWeight_1_weightRead_5_data[1935 : 1928];
  assign dSP_754_b = _zz_b_5[15 : 8];
  assign dSP_755_a = loadWeight_1_weightRead_5_data[1815 : 1808];
  assign dSP_755_d = loadWeight_1_weightRead_5_data[1943 : 1936];
  assign dSP_755_b = _zz_b_5[23 : 16];
  assign dSP_756_a = loadWeight_1_weightRead_5_data[1823 : 1816];
  assign dSP_756_d = loadWeight_1_weightRead_5_data[1951 : 1944];
  assign dSP_756_b = _zz_b_5[31 : 24];
  assign dSP_757_a = loadWeight_1_weightRead_5_data[1831 : 1824];
  assign dSP_757_d = loadWeight_1_weightRead_5_data[1959 : 1952];
  assign dSP_757_b = _zz_b_5[39 : 32];
  assign dSP_758_a = loadWeight_1_weightRead_5_data[1839 : 1832];
  assign dSP_758_d = loadWeight_1_weightRead_5_data[1967 : 1960];
  assign dSP_758_b = _zz_b_5[47 : 40];
  assign dSP_759_a = loadWeight_1_weightRead_5_data[1847 : 1840];
  assign dSP_759_d = loadWeight_1_weightRead_5_data[1975 : 1968];
  assign dSP_759_b = _zz_b_5[55 : 48];
  assign dSP_760_a = loadWeight_1_weightRead_5_data[1855 : 1848];
  assign dSP_760_d = loadWeight_1_weightRead_5_data[1983 : 1976];
  assign dSP_760_b = _zz_b_5[63 : 56];
  assign dSP_761_a = loadWeight_1_weightRead_5_data[1863 : 1856];
  assign dSP_761_d = loadWeight_1_weightRead_5_data[1991 : 1984];
  assign dSP_761_b = _zz_b_5[71 : 64];
  assign dSP_762_a = loadWeight_1_weightRead_5_data[1871 : 1864];
  assign dSP_762_d = loadWeight_1_weightRead_5_data[1999 : 1992];
  assign dSP_762_b = _zz_b_5[79 : 72];
  assign dSP_763_a = loadWeight_1_weightRead_5_data[1879 : 1872];
  assign dSP_763_d = loadWeight_1_weightRead_5_data[2007 : 2000];
  assign dSP_763_b = _zz_b_5[87 : 80];
  assign dSP_764_a = loadWeight_1_weightRead_5_data[1887 : 1880];
  assign dSP_764_d = loadWeight_1_weightRead_5_data[2015 : 2008];
  assign dSP_764_b = _zz_b_5[95 : 88];
  assign dSP_765_a = loadWeight_1_weightRead_5_data[1895 : 1888];
  assign dSP_765_d = loadWeight_1_weightRead_5_data[2023 : 2016];
  assign dSP_765_b = _zz_b_5[103 : 96];
  assign dSP_766_a = loadWeight_1_weightRead_5_data[1903 : 1896];
  assign dSP_766_d = loadWeight_1_weightRead_5_data[2031 : 2024];
  assign dSP_766_b = _zz_b_5[111 : 104];
  assign dSP_767_a = loadWeight_1_weightRead_5_data[1911 : 1904];
  assign dSP_767_d = loadWeight_1_weightRead_5_data[2039 : 2032];
  assign dSP_767_b = _zz_b_5[119 : 112];
  assign dSP_768_a = loadWeight_1_weightRead_5_data[1919 : 1912];
  assign dSP_768_d = loadWeight_1_weightRead_5_data[2047 : 2040];
  assign dSP_768_b = _zz_b_5[127 : 120];
  assign dSP_769_a = loadWeight_1_weightRead_6_data[7 : 0];
  assign dSP_769_d = loadWeight_1_weightRead_6_data[135 : 128];
  assign dSP_769_b = _zz_b_6[7 : 0];
  assign dSP_770_a = loadWeight_1_weightRead_6_data[15 : 8];
  assign dSP_770_d = loadWeight_1_weightRead_6_data[143 : 136];
  assign dSP_770_b = _zz_b_6[15 : 8];
  assign dSP_771_a = loadWeight_1_weightRead_6_data[23 : 16];
  assign dSP_771_d = loadWeight_1_weightRead_6_data[151 : 144];
  assign dSP_771_b = _zz_b_6[23 : 16];
  assign dSP_772_a = loadWeight_1_weightRead_6_data[31 : 24];
  assign dSP_772_d = loadWeight_1_weightRead_6_data[159 : 152];
  assign dSP_772_b = _zz_b_6[31 : 24];
  assign dSP_773_a = loadWeight_1_weightRead_6_data[39 : 32];
  assign dSP_773_d = loadWeight_1_weightRead_6_data[167 : 160];
  assign dSP_773_b = _zz_b_6[39 : 32];
  assign dSP_774_a = loadWeight_1_weightRead_6_data[47 : 40];
  assign dSP_774_d = loadWeight_1_weightRead_6_data[175 : 168];
  assign dSP_774_b = _zz_b_6[47 : 40];
  assign dSP_775_a = loadWeight_1_weightRead_6_data[55 : 48];
  assign dSP_775_d = loadWeight_1_weightRead_6_data[183 : 176];
  assign dSP_775_b = _zz_b_6[55 : 48];
  assign dSP_776_a = loadWeight_1_weightRead_6_data[63 : 56];
  assign dSP_776_d = loadWeight_1_weightRead_6_data[191 : 184];
  assign dSP_776_b = _zz_b_6[63 : 56];
  assign dSP_777_a = loadWeight_1_weightRead_6_data[71 : 64];
  assign dSP_777_d = loadWeight_1_weightRead_6_data[199 : 192];
  assign dSP_777_b = _zz_b_6[71 : 64];
  assign dSP_778_a = loadWeight_1_weightRead_6_data[79 : 72];
  assign dSP_778_d = loadWeight_1_weightRead_6_data[207 : 200];
  assign dSP_778_b = _zz_b_6[79 : 72];
  assign dSP_779_a = loadWeight_1_weightRead_6_data[87 : 80];
  assign dSP_779_d = loadWeight_1_weightRead_6_data[215 : 208];
  assign dSP_779_b = _zz_b_6[87 : 80];
  assign dSP_780_a = loadWeight_1_weightRead_6_data[95 : 88];
  assign dSP_780_d = loadWeight_1_weightRead_6_data[223 : 216];
  assign dSP_780_b = _zz_b_6[95 : 88];
  assign dSP_781_a = loadWeight_1_weightRead_6_data[103 : 96];
  assign dSP_781_d = loadWeight_1_weightRead_6_data[231 : 224];
  assign dSP_781_b = _zz_b_6[103 : 96];
  assign dSP_782_a = loadWeight_1_weightRead_6_data[111 : 104];
  assign dSP_782_d = loadWeight_1_weightRead_6_data[239 : 232];
  assign dSP_782_b = _zz_b_6[111 : 104];
  assign dSP_783_a = loadWeight_1_weightRead_6_data[119 : 112];
  assign dSP_783_d = loadWeight_1_weightRead_6_data[247 : 240];
  assign dSP_783_b = _zz_b_6[119 : 112];
  assign dSP_784_a = loadWeight_1_weightRead_6_data[127 : 120];
  assign dSP_784_d = loadWeight_1_weightRead_6_data[255 : 248];
  assign dSP_784_b = _zz_b_6[127 : 120];
  assign dSP_785_a = loadWeight_1_weightRead_6_data[263 : 256];
  assign dSP_785_d = loadWeight_1_weightRead_6_data[391 : 384];
  assign dSP_785_b = _zz_b_6[7 : 0];
  assign dSP_786_a = loadWeight_1_weightRead_6_data[271 : 264];
  assign dSP_786_d = loadWeight_1_weightRead_6_data[399 : 392];
  assign dSP_786_b = _zz_b_6[15 : 8];
  assign dSP_787_a = loadWeight_1_weightRead_6_data[279 : 272];
  assign dSP_787_d = loadWeight_1_weightRead_6_data[407 : 400];
  assign dSP_787_b = _zz_b_6[23 : 16];
  assign dSP_788_a = loadWeight_1_weightRead_6_data[287 : 280];
  assign dSP_788_d = loadWeight_1_weightRead_6_data[415 : 408];
  assign dSP_788_b = _zz_b_6[31 : 24];
  assign dSP_789_a = loadWeight_1_weightRead_6_data[295 : 288];
  assign dSP_789_d = loadWeight_1_weightRead_6_data[423 : 416];
  assign dSP_789_b = _zz_b_6[39 : 32];
  assign dSP_790_a = loadWeight_1_weightRead_6_data[303 : 296];
  assign dSP_790_d = loadWeight_1_weightRead_6_data[431 : 424];
  assign dSP_790_b = _zz_b_6[47 : 40];
  assign dSP_791_a = loadWeight_1_weightRead_6_data[311 : 304];
  assign dSP_791_d = loadWeight_1_weightRead_6_data[439 : 432];
  assign dSP_791_b = _zz_b_6[55 : 48];
  assign dSP_792_a = loadWeight_1_weightRead_6_data[319 : 312];
  assign dSP_792_d = loadWeight_1_weightRead_6_data[447 : 440];
  assign dSP_792_b = _zz_b_6[63 : 56];
  assign dSP_793_a = loadWeight_1_weightRead_6_data[327 : 320];
  assign dSP_793_d = loadWeight_1_weightRead_6_data[455 : 448];
  assign dSP_793_b = _zz_b_6[71 : 64];
  assign dSP_794_a = loadWeight_1_weightRead_6_data[335 : 328];
  assign dSP_794_d = loadWeight_1_weightRead_6_data[463 : 456];
  assign dSP_794_b = _zz_b_6[79 : 72];
  assign dSP_795_a = loadWeight_1_weightRead_6_data[343 : 336];
  assign dSP_795_d = loadWeight_1_weightRead_6_data[471 : 464];
  assign dSP_795_b = _zz_b_6[87 : 80];
  assign dSP_796_a = loadWeight_1_weightRead_6_data[351 : 344];
  assign dSP_796_d = loadWeight_1_weightRead_6_data[479 : 472];
  assign dSP_796_b = _zz_b_6[95 : 88];
  assign dSP_797_a = loadWeight_1_weightRead_6_data[359 : 352];
  assign dSP_797_d = loadWeight_1_weightRead_6_data[487 : 480];
  assign dSP_797_b = _zz_b_6[103 : 96];
  assign dSP_798_a = loadWeight_1_weightRead_6_data[367 : 360];
  assign dSP_798_d = loadWeight_1_weightRead_6_data[495 : 488];
  assign dSP_798_b = _zz_b_6[111 : 104];
  assign dSP_799_a = loadWeight_1_weightRead_6_data[375 : 368];
  assign dSP_799_d = loadWeight_1_weightRead_6_data[503 : 496];
  assign dSP_799_b = _zz_b_6[119 : 112];
  assign dSP_800_a = loadWeight_1_weightRead_6_data[383 : 376];
  assign dSP_800_d = loadWeight_1_weightRead_6_data[511 : 504];
  assign dSP_800_b = _zz_b_6[127 : 120];
  assign dSP_801_a = loadWeight_1_weightRead_6_data[519 : 512];
  assign dSP_801_d = loadWeight_1_weightRead_6_data[647 : 640];
  assign dSP_801_b = _zz_b_6[7 : 0];
  assign dSP_802_a = loadWeight_1_weightRead_6_data[527 : 520];
  assign dSP_802_d = loadWeight_1_weightRead_6_data[655 : 648];
  assign dSP_802_b = _zz_b_6[15 : 8];
  assign dSP_803_a = loadWeight_1_weightRead_6_data[535 : 528];
  assign dSP_803_d = loadWeight_1_weightRead_6_data[663 : 656];
  assign dSP_803_b = _zz_b_6[23 : 16];
  assign dSP_804_a = loadWeight_1_weightRead_6_data[543 : 536];
  assign dSP_804_d = loadWeight_1_weightRead_6_data[671 : 664];
  assign dSP_804_b = _zz_b_6[31 : 24];
  assign dSP_805_a = loadWeight_1_weightRead_6_data[551 : 544];
  assign dSP_805_d = loadWeight_1_weightRead_6_data[679 : 672];
  assign dSP_805_b = _zz_b_6[39 : 32];
  assign dSP_806_a = loadWeight_1_weightRead_6_data[559 : 552];
  assign dSP_806_d = loadWeight_1_weightRead_6_data[687 : 680];
  assign dSP_806_b = _zz_b_6[47 : 40];
  assign dSP_807_a = loadWeight_1_weightRead_6_data[567 : 560];
  assign dSP_807_d = loadWeight_1_weightRead_6_data[695 : 688];
  assign dSP_807_b = _zz_b_6[55 : 48];
  assign dSP_808_a = loadWeight_1_weightRead_6_data[575 : 568];
  assign dSP_808_d = loadWeight_1_weightRead_6_data[703 : 696];
  assign dSP_808_b = _zz_b_6[63 : 56];
  assign dSP_809_a = loadWeight_1_weightRead_6_data[583 : 576];
  assign dSP_809_d = loadWeight_1_weightRead_6_data[711 : 704];
  assign dSP_809_b = _zz_b_6[71 : 64];
  assign dSP_810_a = loadWeight_1_weightRead_6_data[591 : 584];
  assign dSP_810_d = loadWeight_1_weightRead_6_data[719 : 712];
  assign dSP_810_b = _zz_b_6[79 : 72];
  assign dSP_811_a = loadWeight_1_weightRead_6_data[599 : 592];
  assign dSP_811_d = loadWeight_1_weightRead_6_data[727 : 720];
  assign dSP_811_b = _zz_b_6[87 : 80];
  assign dSP_812_a = loadWeight_1_weightRead_6_data[607 : 600];
  assign dSP_812_d = loadWeight_1_weightRead_6_data[735 : 728];
  assign dSP_812_b = _zz_b_6[95 : 88];
  assign dSP_813_a = loadWeight_1_weightRead_6_data[615 : 608];
  assign dSP_813_d = loadWeight_1_weightRead_6_data[743 : 736];
  assign dSP_813_b = _zz_b_6[103 : 96];
  assign dSP_814_a = loadWeight_1_weightRead_6_data[623 : 616];
  assign dSP_814_d = loadWeight_1_weightRead_6_data[751 : 744];
  assign dSP_814_b = _zz_b_6[111 : 104];
  assign dSP_815_a = loadWeight_1_weightRead_6_data[631 : 624];
  assign dSP_815_d = loadWeight_1_weightRead_6_data[759 : 752];
  assign dSP_815_b = _zz_b_6[119 : 112];
  assign dSP_816_a = loadWeight_1_weightRead_6_data[639 : 632];
  assign dSP_816_d = loadWeight_1_weightRead_6_data[767 : 760];
  assign dSP_816_b = _zz_b_6[127 : 120];
  assign dSP_817_a = loadWeight_1_weightRead_6_data[775 : 768];
  assign dSP_817_d = loadWeight_1_weightRead_6_data[903 : 896];
  assign dSP_817_b = _zz_b_6[7 : 0];
  assign dSP_818_a = loadWeight_1_weightRead_6_data[783 : 776];
  assign dSP_818_d = loadWeight_1_weightRead_6_data[911 : 904];
  assign dSP_818_b = _zz_b_6[15 : 8];
  assign dSP_819_a = loadWeight_1_weightRead_6_data[791 : 784];
  assign dSP_819_d = loadWeight_1_weightRead_6_data[919 : 912];
  assign dSP_819_b = _zz_b_6[23 : 16];
  assign dSP_820_a = loadWeight_1_weightRead_6_data[799 : 792];
  assign dSP_820_d = loadWeight_1_weightRead_6_data[927 : 920];
  assign dSP_820_b = _zz_b_6[31 : 24];
  assign dSP_821_a = loadWeight_1_weightRead_6_data[807 : 800];
  assign dSP_821_d = loadWeight_1_weightRead_6_data[935 : 928];
  assign dSP_821_b = _zz_b_6[39 : 32];
  assign dSP_822_a = loadWeight_1_weightRead_6_data[815 : 808];
  assign dSP_822_d = loadWeight_1_weightRead_6_data[943 : 936];
  assign dSP_822_b = _zz_b_6[47 : 40];
  assign dSP_823_a = loadWeight_1_weightRead_6_data[823 : 816];
  assign dSP_823_d = loadWeight_1_weightRead_6_data[951 : 944];
  assign dSP_823_b = _zz_b_6[55 : 48];
  assign dSP_824_a = loadWeight_1_weightRead_6_data[831 : 824];
  assign dSP_824_d = loadWeight_1_weightRead_6_data[959 : 952];
  assign dSP_824_b = _zz_b_6[63 : 56];
  assign dSP_825_a = loadWeight_1_weightRead_6_data[839 : 832];
  assign dSP_825_d = loadWeight_1_weightRead_6_data[967 : 960];
  assign dSP_825_b = _zz_b_6[71 : 64];
  assign dSP_826_a = loadWeight_1_weightRead_6_data[847 : 840];
  assign dSP_826_d = loadWeight_1_weightRead_6_data[975 : 968];
  assign dSP_826_b = _zz_b_6[79 : 72];
  assign dSP_827_a = loadWeight_1_weightRead_6_data[855 : 848];
  assign dSP_827_d = loadWeight_1_weightRead_6_data[983 : 976];
  assign dSP_827_b = _zz_b_6[87 : 80];
  assign dSP_828_a = loadWeight_1_weightRead_6_data[863 : 856];
  assign dSP_828_d = loadWeight_1_weightRead_6_data[991 : 984];
  assign dSP_828_b = _zz_b_6[95 : 88];
  assign dSP_829_a = loadWeight_1_weightRead_6_data[871 : 864];
  assign dSP_829_d = loadWeight_1_weightRead_6_data[999 : 992];
  assign dSP_829_b = _zz_b_6[103 : 96];
  assign dSP_830_a = loadWeight_1_weightRead_6_data[879 : 872];
  assign dSP_830_d = loadWeight_1_weightRead_6_data[1007 : 1000];
  assign dSP_830_b = _zz_b_6[111 : 104];
  assign dSP_831_a = loadWeight_1_weightRead_6_data[887 : 880];
  assign dSP_831_d = loadWeight_1_weightRead_6_data[1015 : 1008];
  assign dSP_831_b = _zz_b_6[119 : 112];
  assign dSP_832_a = loadWeight_1_weightRead_6_data[895 : 888];
  assign dSP_832_d = loadWeight_1_weightRead_6_data[1023 : 1016];
  assign dSP_832_b = _zz_b_6[127 : 120];
  assign dSP_833_a = loadWeight_1_weightRead_6_data[1031 : 1024];
  assign dSP_833_d = loadWeight_1_weightRead_6_data[1159 : 1152];
  assign dSP_833_b = _zz_b_6[7 : 0];
  assign dSP_834_a = loadWeight_1_weightRead_6_data[1039 : 1032];
  assign dSP_834_d = loadWeight_1_weightRead_6_data[1167 : 1160];
  assign dSP_834_b = _zz_b_6[15 : 8];
  assign dSP_835_a = loadWeight_1_weightRead_6_data[1047 : 1040];
  assign dSP_835_d = loadWeight_1_weightRead_6_data[1175 : 1168];
  assign dSP_835_b = _zz_b_6[23 : 16];
  assign dSP_836_a = loadWeight_1_weightRead_6_data[1055 : 1048];
  assign dSP_836_d = loadWeight_1_weightRead_6_data[1183 : 1176];
  assign dSP_836_b = _zz_b_6[31 : 24];
  assign dSP_837_a = loadWeight_1_weightRead_6_data[1063 : 1056];
  assign dSP_837_d = loadWeight_1_weightRead_6_data[1191 : 1184];
  assign dSP_837_b = _zz_b_6[39 : 32];
  assign dSP_838_a = loadWeight_1_weightRead_6_data[1071 : 1064];
  assign dSP_838_d = loadWeight_1_weightRead_6_data[1199 : 1192];
  assign dSP_838_b = _zz_b_6[47 : 40];
  assign dSP_839_a = loadWeight_1_weightRead_6_data[1079 : 1072];
  assign dSP_839_d = loadWeight_1_weightRead_6_data[1207 : 1200];
  assign dSP_839_b = _zz_b_6[55 : 48];
  assign dSP_840_a = loadWeight_1_weightRead_6_data[1087 : 1080];
  assign dSP_840_d = loadWeight_1_weightRead_6_data[1215 : 1208];
  assign dSP_840_b = _zz_b_6[63 : 56];
  assign dSP_841_a = loadWeight_1_weightRead_6_data[1095 : 1088];
  assign dSP_841_d = loadWeight_1_weightRead_6_data[1223 : 1216];
  assign dSP_841_b = _zz_b_6[71 : 64];
  assign dSP_842_a = loadWeight_1_weightRead_6_data[1103 : 1096];
  assign dSP_842_d = loadWeight_1_weightRead_6_data[1231 : 1224];
  assign dSP_842_b = _zz_b_6[79 : 72];
  assign dSP_843_a = loadWeight_1_weightRead_6_data[1111 : 1104];
  assign dSP_843_d = loadWeight_1_weightRead_6_data[1239 : 1232];
  assign dSP_843_b = _zz_b_6[87 : 80];
  assign dSP_844_a = loadWeight_1_weightRead_6_data[1119 : 1112];
  assign dSP_844_d = loadWeight_1_weightRead_6_data[1247 : 1240];
  assign dSP_844_b = _zz_b_6[95 : 88];
  assign dSP_845_a = loadWeight_1_weightRead_6_data[1127 : 1120];
  assign dSP_845_d = loadWeight_1_weightRead_6_data[1255 : 1248];
  assign dSP_845_b = _zz_b_6[103 : 96];
  assign dSP_846_a = loadWeight_1_weightRead_6_data[1135 : 1128];
  assign dSP_846_d = loadWeight_1_weightRead_6_data[1263 : 1256];
  assign dSP_846_b = _zz_b_6[111 : 104];
  assign dSP_847_a = loadWeight_1_weightRead_6_data[1143 : 1136];
  assign dSP_847_d = loadWeight_1_weightRead_6_data[1271 : 1264];
  assign dSP_847_b = _zz_b_6[119 : 112];
  assign dSP_848_a = loadWeight_1_weightRead_6_data[1151 : 1144];
  assign dSP_848_d = loadWeight_1_weightRead_6_data[1279 : 1272];
  assign dSP_848_b = _zz_b_6[127 : 120];
  assign dSP_849_a = loadWeight_1_weightRead_6_data[1287 : 1280];
  assign dSP_849_d = loadWeight_1_weightRead_6_data[1415 : 1408];
  assign dSP_849_b = _zz_b_6[7 : 0];
  assign dSP_850_a = loadWeight_1_weightRead_6_data[1295 : 1288];
  assign dSP_850_d = loadWeight_1_weightRead_6_data[1423 : 1416];
  assign dSP_850_b = _zz_b_6[15 : 8];
  assign dSP_851_a = loadWeight_1_weightRead_6_data[1303 : 1296];
  assign dSP_851_d = loadWeight_1_weightRead_6_data[1431 : 1424];
  assign dSP_851_b = _zz_b_6[23 : 16];
  assign dSP_852_a = loadWeight_1_weightRead_6_data[1311 : 1304];
  assign dSP_852_d = loadWeight_1_weightRead_6_data[1439 : 1432];
  assign dSP_852_b = _zz_b_6[31 : 24];
  assign dSP_853_a = loadWeight_1_weightRead_6_data[1319 : 1312];
  assign dSP_853_d = loadWeight_1_weightRead_6_data[1447 : 1440];
  assign dSP_853_b = _zz_b_6[39 : 32];
  assign dSP_854_a = loadWeight_1_weightRead_6_data[1327 : 1320];
  assign dSP_854_d = loadWeight_1_weightRead_6_data[1455 : 1448];
  assign dSP_854_b = _zz_b_6[47 : 40];
  assign dSP_855_a = loadWeight_1_weightRead_6_data[1335 : 1328];
  assign dSP_855_d = loadWeight_1_weightRead_6_data[1463 : 1456];
  assign dSP_855_b = _zz_b_6[55 : 48];
  assign dSP_856_a = loadWeight_1_weightRead_6_data[1343 : 1336];
  assign dSP_856_d = loadWeight_1_weightRead_6_data[1471 : 1464];
  assign dSP_856_b = _zz_b_6[63 : 56];
  assign dSP_857_a = loadWeight_1_weightRead_6_data[1351 : 1344];
  assign dSP_857_d = loadWeight_1_weightRead_6_data[1479 : 1472];
  assign dSP_857_b = _zz_b_6[71 : 64];
  assign dSP_858_a = loadWeight_1_weightRead_6_data[1359 : 1352];
  assign dSP_858_d = loadWeight_1_weightRead_6_data[1487 : 1480];
  assign dSP_858_b = _zz_b_6[79 : 72];
  assign dSP_859_a = loadWeight_1_weightRead_6_data[1367 : 1360];
  assign dSP_859_d = loadWeight_1_weightRead_6_data[1495 : 1488];
  assign dSP_859_b = _zz_b_6[87 : 80];
  assign dSP_860_a = loadWeight_1_weightRead_6_data[1375 : 1368];
  assign dSP_860_d = loadWeight_1_weightRead_6_data[1503 : 1496];
  assign dSP_860_b = _zz_b_6[95 : 88];
  assign dSP_861_a = loadWeight_1_weightRead_6_data[1383 : 1376];
  assign dSP_861_d = loadWeight_1_weightRead_6_data[1511 : 1504];
  assign dSP_861_b = _zz_b_6[103 : 96];
  assign dSP_862_a = loadWeight_1_weightRead_6_data[1391 : 1384];
  assign dSP_862_d = loadWeight_1_weightRead_6_data[1519 : 1512];
  assign dSP_862_b = _zz_b_6[111 : 104];
  assign dSP_863_a = loadWeight_1_weightRead_6_data[1399 : 1392];
  assign dSP_863_d = loadWeight_1_weightRead_6_data[1527 : 1520];
  assign dSP_863_b = _zz_b_6[119 : 112];
  assign dSP_864_a = loadWeight_1_weightRead_6_data[1407 : 1400];
  assign dSP_864_d = loadWeight_1_weightRead_6_data[1535 : 1528];
  assign dSP_864_b = _zz_b_6[127 : 120];
  assign dSP_865_a = loadWeight_1_weightRead_6_data[1543 : 1536];
  assign dSP_865_d = loadWeight_1_weightRead_6_data[1671 : 1664];
  assign dSP_865_b = _zz_b_6[7 : 0];
  assign dSP_866_a = loadWeight_1_weightRead_6_data[1551 : 1544];
  assign dSP_866_d = loadWeight_1_weightRead_6_data[1679 : 1672];
  assign dSP_866_b = _zz_b_6[15 : 8];
  assign dSP_867_a = loadWeight_1_weightRead_6_data[1559 : 1552];
  assign dSP_867_d = loadWeight_1_weightRead_6_data[1687 : 1680];
  assign dSP_867_b = _zz_b_6[23 : 16];
  assign dSP_868_a = loadWeight_1_weightRead_6_data[1567 : 1560];
  assign dSP_868_d = loadWeight_1_weightRead_6_data[1695 : 1688];
  assign dSP_868_b = _zz_b_6[31 : 24];
  assign dSP_869_a = loadWeight_1_weightRead_6_data[1575 : 1568];
  assign dSP_869_d = loadWeight_1_weightRead_6_data[1703 : 1696];
  assign dSP_869_b = _zz_b_6[39 : 32];
  assign dSP_870_a = loadWeight_1_weightRead_6_data[1583 : 1576];
  assign dSP_870_d = loadWeight_1_weightRead_6_data[1711 : 1704];
  assign dSP_870_b = _zz_b_6[47 : 40];
  assign dSP_871_a = loadWeight_1_weightRead_6_data[1591 : 1584];
  assign dSP_871_d = loadWeight_1_weightRead_6_data[1719 : 1712];
  assign dSP_871_b = _zz_b_6[55 : 48];
  assign dSP_872_a = loadWeight_1_weightRead_6_data[1599 : 1592];
  assign dSP_872_d = loadWeight_1_weightRead_6_data[1727 : 1720];
  assign dSP_872_b = _zz_b_6[63 : 56];
  assign dSP_873_a = loadWeight_1_weightRead_6_data[1607 : 1600];
  assign dSP_873_d = loadWeight_1_weightRead_6_data[1735 : 1728];
  assign dSP_873_b = _zz_b_6[71 : 64];
  assign dSP_874_a = loadWeight_1_weightRead_6_data[1615 : 1608];
  assign dSP_874_d = loadWeight_1_weightRead_6_data[1743 : 1736];
  assign dSP_874_b = _zz_b_6[79 : 72];
  assign dSP_875_a = loadWeight_1_weightRead_6_data[1623 : 1616];
  assign dSP_875_d = loadWeight_1_weightRead_6_data[1751 : 1744];
  assign dSP_875_b = _zz_b_6[87 : 80];
  assign dSP_876_a = loadWeight_1_weightRead_6_data[1631 : 1624];
  assign dSP_876_d = loadWeight_1_weightRead_6_data[1759 : 1752];
  assign dSP_876_b = _zz_b_6[95 : 88];
  assign dSP_877_a = loadWeight_1_weightRead_6_data[1639 : 1632];
  assign dSP_877_d = loadWeight_1_weightRead_6_data[1767 : 1760];
  assign dSP_877_b = _zz_b_6[103 : 96];
  assign dSP_878_a = loadWeight_1_weightRead_6_data[1647 : 1640];
  assign dSP_878_d = loadWeight_1_weightRead_6_data[1775 : 1768];
  assign dSP_878_b = _zz_b_6[111 : 104];
  assign dSP_879_a = loadWeight_1_weightRead_6_data[1655 : 1648];
  assign dSP_879_d = loadWeight_1_weightRead_6_data[1783 : 1776];
  assign dSP_879_b = _zz_b_6[119 : 112];
  assign dSP_880_a = loadWeight_1_weightRead_6_data[1663 : 1656];
  assign dSP_880_d = loadWeight_1_weightRead_6_data[1791 : 1784];
  assign dSP_880_b = _zz_b_6[127 : 120];
  assign dSP_881_a = loadWeight_1_weightRead_6_data[1799 : 1792];
  assign dSP_881_d = loadWeight_1_weightRead_6_data[1927 : 1920];
  assign dSP_881_b = _zz_b_6[7 : 0];
  assign dSP_882_a = loadWeight_1_weightRead_6_data[1807 : 1800];
  assign dSP_882_d = loadWeight_1_weightRead_6_data[1935 : 1928];
  assign dSP_882_b = _zz_b_6[15 : 8];
  assign dSP_883_a = loadWeight_1_weightRead_6_data[1815 : 1808];
  assign dSP_883_d = loadWeight_1_weightRead_6_data[1943 : 1936];
  assign dSP_883_b = _zz_b_6[23 : 16];
  assign dSP_884_a = loadWeight_1_weightRead_6_data[1823 : 1816];
  assign dSP_884_d = loadWeight_1_weightRead_6_data[1951 : 1944];
  assign dSP_884_b = _zz_b_6[31 : 24];
  assign dSP_885_a = loadWeight_1_weightRead_6_data[1831 : 1824];
  assign dSP_885_d = loadWeight_1_weightRead_6_data[1959 : 1952];
  assign dSP_885_b = _zz_b_6[39 : 32];
  assign dSP_886_a = loadWeight_1_weightRead_6_data[1839 : 1832];
  assign dSP_886_d = loadWeight_1_weightRead_6_data[1967 : 1960];
  assign dSP_886_b = _zz_b_6[47 : 40];
  assign dSP_887_a = loadWeight_1_weightRead_6_data[1847 : 1840];
  assign dSP_887_d = loadWeight_1_weightRead_6_data[1975 : 1968];
  assign dSP_887_b = _zz_b_6[55 : 48];
  assign dSP_888_a = loadWeight_1_weightRead_6_data[1855 : 1848];
  assign dSP_888_d = loadWeight_1_weightRead_6_data[1983 : 1976];
  assign dSP_888_b = _zz_b_6[63 : 56];
  assign dSP_889_a = loadWeight_1_weightRead_6_data[1863 : 1856];
  assign dSP_889_d = loadWeight_1_weightRead_6_data[1991 : 1984];
  assign dSP_889_b = _zz_b_6[71 : 64];
  assign dSP_890_a = loadWeight_1_weightRead_6_data[1871 : 1864];
  assign dSP_890_d = loadWeight_1_weightRead_6_data[1999 : 1992];
  assign dSP_890_b = _zz_b_6[79 : 72];
  assign dSP_891_a = loadWeight_1_weightRead_6_data[1879 : 1872];
  assign dSP_891_d = loadWeight_1_weightRead_6_data[2007 : 2000];
  assign dSP_891_b = _zz_b_6[87 : 80];
  assign dSP_892_a = loadWeight_1_weightRead_6_data[1887 : 1880];
  assign dSP_892_d = loadWeight_1_weightRead_6_data[2015 : 2008];
  assign dSP_892_b = _zz_b_6[95 : 88];
  assign dSP_893_a = loadWeight_1_weightRead_6_data[1895 : 1888];
  assign dSP_893_d = loadWeight_1_weightRead_6_data[2023 : 2016];
  assign dSP_893_b = _zz_b_6[103 : 96];
  assign dSP_894_a = loadWeight_1_weightRead_6_data[1903 : 1896];
  assign dSP_894_d = loadWeight_1_weightRead_6_data[2031 : 2024];
  assign dSP_894_b = _zz_b_6[111 : 104];
  assign dSP_895_a = loadWeight_1_weightRead_6_data[1911 : 1904];
  assign dSP_895_d = loadWeight_1_weightRead_6_data[2039 : 2032];
  assign dSP_895_b = _zz_b_6[119 : 112];
  assign dSP_896_a = loadWeight_1_weightRead_6_data[1919 : 1912];
  assign dSP_896_d = loadWeight_1_weightRead_6_data[2047 : 2040];
  assign dSP_896_b = _zz_b_6[127 : 120];
  assign dSP_897_a = loadWeight_1_weightRead_7_data[7 : 0];
  assign dSP_897_d = loadWeight_1_weightRead_7_data[135 : 128];
  assign dSP_897_b = _zz_b_7[7 : 0];
  assign dSP_898_a = loadWeight_1_weightRead_7_data[15 : 8];
  assign dSP_898_d = loadWeight_1_weightRead_7_data[143 : 136];
  assign dSP_898_b = _zz_b_7[15 : 8];
  assign dSP_899_a = loadWeight_1_weightRead_7_data[23 : 16];
  assign dSP_899_d = loadWeight_1_weightRead_7_data[151 : 144];
  assign dSP_899_b = _zz_b_7[23 : 16];
  assign dSP_900_a = loadWeight_1_weightRead_7_data[31 : 24];
  assign dSP_900_d = loadWeight_1_weightRead_7_data[159 : 152];
  assign dSP_900_b = _zz_b_7[31 : 24];
  assign dSP_901_a = loadWeight_1_weightRead_7_data[39 : 32];
  assign dSP_901_d = loadWeight_1_weightRead_7_data[167 : 160];
  assign dSP_901_b = _zz_b_7[39 : 32];
  assign dSP_902_a = loadWeight_1_weightRead_7_data[47 : 40];
  assign dSP_902_d = loadWeight_1_weightRead_7_data[175 : 168];
  assign dSP_902_b = _zz_b_7[47 : 40];
  assign dSP_903_a = loadWeight_1_weightRead_7_data[55 : 48];
  assign dSP_903_d = loadWeight_1_weightRead_7_data[183 : 176];
  assign dSP_903_b = _zz_b_7[55 : 48];
  assign dSP_904_a = loadWeight_1_weightRead_7_data[63 : 56];
  assign dSP_904_d = loadWeight_1_weightRead_7_data[191 : 184];
  assign dSP_904_b = _zz_b_7[63 : 56];
  assign dSP_905_a = loadWeight_1_weightRead_7_data[71 : 64];
  assign dSP_905_d = loadWeight_1_weightRead_7_data[199 : 192];
  assign dSP_905_b = _zz_b_7[71 : 64];
  assign dSP_906_a = loadWeight_1_weightRead_7_data[79 : 72];
  assign dSP_906_d = loadWeight_1_weightRead_7_data[207 : 200];
  assign dSP_906_b = _zz_b_7[79 : 72];
  assign dSP_907_a = loadWeight_1_weightRead_7_data[87 : 80];
  assign dSP_907_d = loadWeight_1_weightRead_7_data[215 : 208];
  assign dSP_907_b = _zz_b_7[87 : 80];
  assign dSP_908_a = loadWeight_1_weightRead_7_data[95 : 88];
  assign dSP_908_d = loadWeight_1_weightRead_7_data[223 : 216];
  assign dSP_908_b = _zz_b_7[95 : 88];
  assign dSP_909_a = loadWeight_1_weightRead_7_data[103 : 96];
  assign dSP_909_d = loadWeight_1_weightRead_7_data[231 : 224];
  assign dSP_909_b = _zz_b_7[103 : 96];
  assign dSP_910_a = loadWeight_1_weightRead_7_data[111 : 104];
  assign dSP_910_d = loadWeight_1_weightRead_7_data[239 : 232];
  assign dSP_910_b = _zz_b_7[111 : 104];
  assign dSP_911_a = loadWeight_1_weightRead_7_data[119 : 112];
  assign dSP_911_d = loadWeight_1_weightRead_7_data[247 : 240];
  assign dSP_911_b = _zz_b_7[119 : 112];
  assign dSP_912_a = loadWeight_1_weightRead_7_data[127 : 120];
  assign dSP_912_d = loadWeight_1_weightRead_7_data[255 : 248];
  assign dSP_912_b = _zz_b_7[127 : 120];
  assign dSP_913_a = loadWeight_1_weightRead_7_data[263 : 256];
  assign dSP_913_d = loadWeight_1_weightRead_7_data[391 : 384];
  assign dSP_913_b = _zz_b_7[7 : 0];
  assign dSP_914_a = loadWeight_1_weightRead_7_data[271 : 264];
  assign dSP_914_d = loadWeight_1_weightRead_7_data[399 : 392];
  assign dSP_914_b = _zz_b_7[15 : 8];
  assign dSP_915_a = loadWeight_1_weightRead_7_data[279 : 272];
  assign dSP_915_d = loadWeight_1_weightRead_7_data[407 : 400];
  assign dSP_915_b = _zz_b_7[23 : 16];
  assign dSP_916_a = loadWeight_1_weightRead_7_data[287 : 280];
  assign dSP_916_d = loadWeight_1_weightRead_7_data[415 : 408];
  assign dSP_916_b = _zz_b_7[31 : 24];
  assign dSP_917_a = loadWeight_1_weightRead_7_data[295 : 288];
  assign dSP_917_d = loadWeight_1_weightRead_7_data[423 : 416];
  assign dSP_917_b = _zz_b_7[39 : 32];
  assign dSP_918_a = loadWeight_1_weightRead_7_data[303 : 296];
  assign dSP_918_d = loadWeight_1_weightRead_7_data[431 : 424];
  assign dSP_918_b = _zz_b_7[47 : 40];
  assign dSP_919_a = loadWeight_1_weightRead_7_data[311 : 304];
  assign dSP_919_d = loadWeight_1_weightRead_7_data[439 : 432];
  assign dSP_919_b = _zz_b_7[55 : 48];
  assign dSP_920_a = loadWeight_1_weightRead_7_data[319 : 312];
  assign dSP_920_d = loadWeight_1_weightRead_7_data[447 : 440];
  assign dSP_920_b = _zz_b_7[63 : 56];
  assign dSP_921_a = loadWeight_1_weightRead_7_data[327 : 320];
  assign dSP_921_d = loadWeight_1_weightRead_7_data[455 : 448];
  assign dSP_921_b = _zz_b_7[71 : 64];
  assign dSP_922_a = loadWeight_1_weightRead_7_data[335 : 328];
  assign dSP_922_d = loadWeight_1_weightRead_7_data[463 : 456];
  assign dSP_922_b = _zz_b_7[79 : 72];
  assign dSP_923_a = loadWeight_1_weightRead_7_data[343 : 336];
  assign dSP_923_d = loadWeight_1_weightRead_7_data[471 : 464];
  assign dSP_923_b = _zz_b_7[87 : 80];
  assign dSP_924_a = loadWeight_1_weightRead_7_data[351 : 344];
  assign dSP_924_d = loadWeight_1_weightRead_7_data[479 : 472];
  assign dSP_924_b = _zz_b_7[95 : 88];
  assign dSP_925_a = loadWeight_1_weightRead_7_data[359 : 352];
  assign dSP_925_d = loadWeight_1_weightRead_7_data[487 : 480];
  assign dSP_925_b = _zz_b_7[103 : 96];
  assign dSP_926_a = loadWeight_1_weightRead_7_data[367 : 360];
  assign dSP_926_d = loadWeight_1_weightRead_7_data[495 : 488];
  assign dSP_926_b = _zz_b_7[111 : 104];
  assign dSP_927_a = loadWeight_1_weightRead_7_data[375 : 368];
  assign dSP_927_d = loadWeight_1_weightRead_7_data[503 : 496];
  assign dSP_927_b = _zz_b_7[119 : 112];
  assign dSP_928_a = loadWeight_1_weightRead_7_data[383 : 376];
  assign dSP_928_d = loadWeight_1_weightRead_7_data[511 : 504];
  assign dSP_928_b = _zz_b_7[127 : 120];
  assign dSP_929_a = loadWeight_1_weightRead_7_data[519 : 512];
  assign dSP_929_d = loadWeight_1_weightRead_7_data[647 : 640];
  assign dSP_929_b = _zz_b_7[7 : 0];
  assign dSP_930_a = loadWeight_1_weightRead_7_data[527 : 520];
  assign dSP_930_d = loadWeight_1_weightRead_7_data[655 : 648];
  assign dSP_930_b = _zz_b_7[15 : 8];
  assign dSP_931_a = loadWeight_1_weightRead_7_data[535 : 528];
  assign dSP_931_d = loadWeight_1_weightRead_7_data[663 : 656];
  assign dSP_931_b = _zz_b_7[23 : 16];
  assign dSP_932_a = loadWeight_1_weightRead_7_data[543 : 536];
  assign dSP_932_d = loadWeight_1_weightRead_7_data[671 : 664];
  assign dSP_932_b = _zz_b_7[31 : 24];
  assign dSP_933_a = loadWeight_1_weightRead_7_data[551 : 544];
  assign dSP_933_d = loadWeight_1_weightRead_7_data[679 : 672];
  assign dSP_933_b = _zz_b_7[39 : 32];
  assign dSP_934_a = loadWeight_1_weightRead_7_data[559 : 552];
  assign dSP_934_d = loadWeight_1_weightRead_7_data[687 : 680];
  assign dSP_934_b = _zz_b_7[47 : 40];
  assign dSP_935_a = loadWeight_1_weightRead_7_data[567 : 560];
  assign dSP_935_d = loadWeight_1_weightRead_7_data[695 : 688];
  assign dSP_935_b = _zz_b_7[55 : 48];
  assign dSP_936_a = loadWeight_1_weightRead_7_data[575 : 568];
  assign dSP_936_d = loadWeight_1_weightRead_7_data[703 : 696];
  assign dSP_936_b = _zz_b_7[63 : 56];
  assign dSP_937_a = loadWeight_1_weightRead_7_data[583 : 576];
  assign dSP_937_d = loadWeight_1_weightRead_7_data[711 : 704];
  assign dSP_937_b = _zz_b_7[71 : 64];
  assign dSP_938_a = loadWeight_1_weightRead_7_data[591 : 584];
  assign dSP_938_d = loadWeight_1_weightRead_7_data[719 : 712];
  assign dSP_938_b = _zz_b_7[79 : 72];
  assign dSP_939_a = loadWeight_1_weightRead_7_data[599 : 592];
  assign dSP_939_d = loadWeight_1_weightRead_7_data[727 : 720];
  assign dSP_939_b = _zz_b_7[87 : 80];
  assign dSP_940_a = loadWeight_1_weightRead_7_data[607 : 600];
  assign dSP_940_d = loadWeight_1_weightRead_7_data[735 : 728];
  assign dSP_940_b = _zz_b_7[95 : 88];
  assign dSP_941_a = loadWeight_1_weightRead_7_data[615 : 608];
  assign dSP_941_d = loadWeight_1_weightRead_7_data[743 : 736];
  assign dSP_941_b = _zz_b_7[103 : 96];
  assign dSP_942_a = loadWeight_1_weightRead_7_data[623 : 616];
  assign dSP_942_d = loadWeight_1_weightRead_7_data[751 : 744];
  assign dSP_942_b = _zz_b_7[111 : 104];
  assign dSP_943_a = loadWeight_1_weightRead_7_data[631 : 624];
  assign dSP_943_d = loadWeight_1_weightRead_7_data[759 : 752];
  assign dSP_943_b = _zz_b_7[119 : 112];
  assign dSP_944_a = loadWeight_1_weightRead_7_data[639 : 632];
  assign dSP_944_d = loadWeight_1_weightRead_7_data[767 : 760];
  assign dSP_944_b = _zz_b_7[127 : 120];
  assign dSP_945_a = loadWeight_1_weightRead_7_data[775 : 768];
  assign dSP_945_d = loadWeight_1_weightRead_7_data[903 : 896];
  assign dSP_945_b = _zz_b_7[7 : 0];
  assign dSP_946_a = loadWeight_1_weightRead_7_data[783 : 776];
  assign dSP_946_d = loadWeight_1_weightRead_7_data[911 : 904];
  assign dSP_946_b = _zz_b_7[15 : 8];
  assign dSP_947_a = loadWeight_1_weightRead_7_data[791 : 784];
  assign dSP_947_d = loadWeight_1_weightRead_7_data[919 : 912];
  assign dSP_947_b = _zz_b_7[23 : 16];
  assign dSP_948_a = loadWeight_1_weightRead_7_data[799 : 792];
  assign dSP_948_d = loadWeight_1_weightRead_7_data[927 : 920];
  assign dSP_948_b = _zz_b_7[31 : 24];
  assign dSP_949_a = loadWeight_1_weightRead_7_data[807 : 800];
  assign dSP_949_d = loadWeight_1_weightRead_7_data[935 : 928];
  assign dSP_949_b = _zz_b_7[39 : 32];
  assign dSP_950_a = loadWeight_1_weightRead_7_data[815 : 808];
  assign dSP_950_d = loadWeight_1_weightRead_7_data[943 : 936];
  assign dSP_950_b = _zz_b_7[47 : 40];
  assign dSP_951_a = loadWeight_1_weightRead_7_data[823 : 816];
  assign dSP_951_d = loadWeight_1_weightRead_7_data[951 : 944];
  assign dSP_951_b = _zz_b_7[55 : 48];
  assign dSP_952_a = loadWeight_1_weightRead_7_data[831 : 824];
  assign dSP_952_d = loadWeight_1_weightRead_7_data[959 : 952];
  assign dSP_952_b = _zz_b_7[63 : 56];
  assign dSP_953_a = loadWeight_1_weightRead_7_data[839 : 832];
  assign dSP_953_d = loadWeight_1_weightRead_7_data[967 : 960];
  assign dSP_953_b = _zz_b_7[71 : 64];
  assign dSP_954_a = loadWeight_1_weightRead_7_data[847 : 840];
  assign dSP_954_d = loadWeight_1_weightRead_7_data[975 : 968];
  assign dSP_954_b = _zz_b_7[79 : 72];
  assign dSP_955_a = loadWeight_1_weightRead_7_data[855 : 848];
  assign dSP_955_d = loadWeight_1_weightRead_7_data[983 : 976];
  assign dSP_955_b = _zz_b_7[87 : 80];
  assign dSP_956_a = loadWeight_1_weightRead_7_data[863 : 856];
  assign dSP_956_d = loadWeight_1_weightRead_7_data[991 : 984];
  assign dSP_956_b = _zz_b_7[95 : 88];
  assign dSP_957_a = loadWeight_1_weightRead_7_data[871 : 864];
  assign dSP_957_d = loadWeight_1_weightRead_7_data[999 : 992];
  assign dSP_957_b = _zz_b_7[103 : 96];
  assign dSP_958_a = loadWeight_1_weightRead_7_data[879 : 872];
  assign dSP_958_d = loadWeight_1_weightRead_7_data[1007 : 1000];
  assign dSP_958_b = _zz_b_7[111 : 104];
  assign dSP_959_a = loadWeight_1_weightRead_7_data[887 : 880];
  assign dSP_959_d = loadWeight_1_weightRead_7_data[1015 : 1008];
  assign dSP_959_b = _zz_b_7[119 : 112];
  assign dSP_960_a = loadWeight_1_weightRead_7_data[895 : 888];
  assign dSP_960_d = loadWeight_1_weightRead_7_data[1023 : 1016];
  assign dSP_960_b = _zz_b_7[127 : 120];
  assign dSP_961_a = loadWeight_1_weightRead_7_data[1031 : 1024];
  assign dSP_961_d = loadWeight_1_weightRead_7_data[1159 : 1152];
  assign dSP_961_b = _zz_b_7[7 : 0];
  assign dSP_962_a = loadWeight_1_weightRead_7_data[1039 : 1032];
  assign dSP_962_d = loadWeight_1_weightRead_7_data[1167 : 1160];
  assign dSP_962_b = _zz_b_7[15 : 8];
  assign dSP_963_a = loadWeight_1_weightRead_7_data[1047 : 1040];
  assign dSP_963_d = loadWeight_1_weightRead_7_data[1175 : 1168];
  assign dSP_963_b = _zz_b_7[23 : 16];
  assign dSP_964_a = loadWeight_1_weightRead_7_data[1055 : 1048];
  assign dSP_964_d = loadWeight_1_weightRead_7_data[1183 : 1176];
  assign dSP_964_b = _zz_b_7[31 : 24];
  assign dSP_965_a = loadWeight_1_weightRead_7_data[1063 : 1056];
  assign dSP_965_d = loadWeight_1_weightRead_7_data[1191 : 1184];
  assign dSP_965_b = _zz_b_7[39 : 32];
  assign dSP_966_a = loadWeight_1_weightRead_7_data[1071 : 1064];
  assign dSP_966_d = loadWeight_1_weightRead_7_data[1199 : 1192];
  assign dSP_966_b = _zz_b_7[47 : 40];
  assign dSP_967_a = loadWeight_1_weightRead_7_data[1079 : 1072];
  assign dSP_967_d = loadWeight_1_weightRead_7_data[1207 : 1200];
  assign dSP_967_b = _zz_b_7[55 : 48];
  assign dSP_968_a = loadWeight_1_weightRead_7_data[1087 : 1080];
  assign dSP_968_d = loadWeight_1_weightRead_7_data[1215 : 1208];
  assign dSP_968_b = _zz_b_7[63 : 56];
  assign dSP_969_a = loadWeight_1_weightRead_7_data[1095 : 1088];
  assign dSP_969_d = loadWeight_1_weightRead_7_data[1223 : 1216];
  assign dSP_969_b = _zz_b_7[71 : 64];
  assign dSP_970_a = loadWeight_1_weightRead_7_data[1103 : 1096];
  assign dSP_970_d = loadWeight_1_weightRead_7_data[1231 : 1224];
  assign dSP_970_b = _zz_b_7[79 : 72];
  assign dSP_971_a = loadWeight_1_weightRead_7_data[1111 : 1104];
  assign dSP_971_d = loadWeight_1_weightRead_7_data[1239 : 1232];
  assign dSP_971_b = _zz_b_7[87 : 80];
  assign dSP_972_a = loadWeight_1_weightRead_7_data[1119 : 1112];
  assign dSP_972_d = loadWeight_1_weightRead_7_data[1247 : 1240];
  assign dSP_972_b = _zz_b_7[95 : 88];
  assign dSP_973_a = loadWeight_1_weightRead_7_data[1127 : 1120];
  assign dSP_973_d = loadWeight_1_weightRead_7_data[1255 : 1248];
  assign dSP_973_b = _zz_b_7[103 : 96];
  assign dSP_974_a = loadWeight_1_weightRead_7_data[1135 : 1128];
  assign dSP_974_d = loadWeight_1_weightRead_7_data[1263 : 1256];
  assign dSP_974_b = _zz_b_7[111 : 104];
  assign dSP_975_a = loadWeight_1_weightRead_7_data[1143 : 1136];
  assign dSP_975_d = loadWeight_1_weightRead_7_data[1271 : 1264];
  assign dSP_975_b = _zz_b_7[119 : 112];
  assign dSP_976_a = loadWeight_1_weightRead_7_data[1151 : 1144];
  assign dSP_976_d = loadWeight_1_weightRead_7_data[1279 : 1272];
  assign dSP_976_b = _zz_b_7[127 : 120];
  assign dSP_977_a = loadWeight_1_weightRead_7_data[1287 : 1280];
  assign dSP_977_d = loadWeight_1_weightRead_7_data[1415 : 1408];
  assign dSP_977_b = _zz_b_7[7 : 0];
  assign dSP_978_a = loadWeight_1_weightRead_7_data[1295 : 1288];
  assign dSP_978_d = loadWeight_1_weightRead_7_data[1423 : 1416];
  assign dSP_978_b = _zz_b_7[15 : 8];
  assign dSP_979_a = loadWeight_1_weightRead_7_data[1303 : 1296];
  assign dSP_979_d = loadWeight_1_weightRead_7_data[1431 : 1424];
  assign dSP_979_b = _zz_b_7[23 : 16];
  assign dSP_980_a = loadWeight_1_weightRead_7_data[1311 : 1304];
  assign dSP_980_d = loadWeight_1_weightRead_7_data[1439 : 1432];
  assign dSP_980_b = _zz_b_7[31 : 24];
  assign dSP_981_a = loadWeight_1_weightRead_7_data[1319 : 1312];
  assign dSP_981_d = loadWeight_1_weightRead_7_data[1447 : 1440];
  assign dSP_981_b = _zz_b_7[39 : 32];
  assign dSP_982_a = loadWeight_1_weightRead_7_data[1327 : 1320];
  assign dSP_982_d = loadWeight_1_weightRead_7_data[1455 : 1448];
  assign dSP_982_b = _zz_b_7[47 : 40];
  assign dSP_983_a = loadWeight_1_weightRead_7_data[1335 : 1328];
  assign dSP_983_d = loadWeight_1_weightRead_7_data[1463 : 1456];
  assign dSP_983_b = _zz_b_7[55 : 48];
  assign dSP_984_a = loadWeight_1_weightRead_7_data[1343 : 1336];
  assign dSP_984_d = loadWeight_1_weightRead_7_data[1471 : 1464];
  assign dSP_984_b = _zz_b_7[63 : 56];
  assign dSP_985_a = loadWeight_1_weightRead_7_data[1351 : 1344];
  assign dSP_985_d = loadWeight_1_weightRead_7_data[1479 : 1472];
  assign dSP_985_b = _zz_b_7[71 : 64];
  assign dSP_986_a = loadWeight_1_weightRead_7_data[1359 : 1352];
  assign dSP_986_d = loadWeight_1_weightRead_7_data[1487 : 1480];
  assign dSP_986_b = _zz_b_7[79 : 72];
  assign dSP_987_a = loadWeight_1_weightRead_7_data[1367 : 1360];
  assign dSP_987_d = loadWeight_1_weightRead_7_data[1495 : 1488];
  assign dSP_987_b = _zz_b_7[87 : 80];
  assign dSP_988_a = loadWeight_1_weightRead_7_data[1375 : 1368];
  assign dSP_988_d = loadWeight_1_weightRead_7_data[1503 : 1496];
  assign dSP_988_b = _zz_b_7[95 : 88];
  assign dSP_989_a = loadWeight_1_weightRead_7_data[1383 : 1376];
  assign dSP_989_d = loadWeight_1_weightRead_7_data[1511 : 1504];
  assign dSP_989_b = _zz_b_7[103 : 96];
  assign dSP_990_a = loadWeight_1_weightRead_7_data[1391 : 1384];
  assign dSP_990_d = loadWeight_1_weightRead_7_data[1519 : 1512];
  assign dSP_990_b = _zz_b_7[111 : 104];
  assign dSP_991_a = loadWeight_1_weightRead_7_data[1399 : 1392];
  assign dSP_991_d = loadWeight_1_weightRead_7_data[1527 : 1520];
  assign dSP_991_b = _zz_b_7[119 : 112];
  assign dSP_992_a = loadWeight_1_weightRead_7_data[1407 : 1400];
  assign dSP_992_d = loadWeight_1_weightRead_7_data[1535 : 1528];
  assign dSP_992_b = _zz_b_7[127 : 120];
  assign dSP_993_a = loadWeight_1_weightRead_7_data[1543 : 1536];
  assign dSP_993_d = loadWeight_1_weightRead_7_data[1671 : 1664];
  assign dSP_993_b = _zz_b_7[7 : 0];
  assign dSP_994_a = loadWeight_1_weightRead_7_data[1551 : 1544];
  assign dSP_994_d = loadWeight_1_weightRead_7_data[1679 : 1672];
  assign dSP_994_b = _zz_b_7[15 : 8];
  assign dSP_995_a = loadWeight_1_weightRead_7_data[1559 : 1552];
  assign dSP_995_d = loadWeight_1_weightRead_7_data[1687 : 1680];
  assign dSP_995_b = _zz_b_7[23 : 16];
  assign dSP_996_a = loadWeight_1_weightRead_7_data[1567 : 1560];
  assign dSP_996_d = loadWeight_1_weightRead_7_data[1695 : 1688];
  assign dSP_996_b = _zz_b_7[31 : 24];
  assign dSP_997_a = loadWeight_1_weightRead_7_data[1575 : 1568];
  assign dSP_997_d = loadWeight_1_weightRead_7_data[1703 : 1696];
  assign dSP_997_b = _zz_b_7[39 : 32];
  assign dSP_998_a = loadWeight_1_weightRead_7_data[1583 : 1576];
  assign dSP_998_d = loadWeight_1_weightRead_7_data[1711 : 1704];
  assign dSP_998_b = _zz_b_7[47 : 40];
  assign dSP_999_a = loadWeight_1_weightRead_7_data[1591 : 1584];
  assign dSP_999_d = loadWeight_1_weightRead_7_data[1719 : 1712];
  assign dSP_999_b = _zz_b_7[55 : 48];
  assign dSP_1000_a = loadWeight_1_weightRead_7_data[1599 : 1592];
  assign dSP_1000_d = loadWeight_1_weightRead_7_data[1727 : 1720];
  assign dSP_1000_b = _zz_b_7[63 : 56];
  assign dSP_1001_a = loadWeight_1_weightRead_7_data[1607 : 1600];
  assign dSP_1001_d = loadWeight_1_weightRead_7_data[1735 : 1728];
  assign dSP_1001_b = _zz_b_7[71 : 64];
  assign dSP_1002_a = loadWeight_1_weightRead_7_data[1615 : 1608];
  assign dSP_1002_d = loadWeight_1_weightRead_7_data[1743 : 1736];
  assign dSP_1002_b = _zz_b_7[79 : 72];
  assign dSP_1003_a = loadWeight_1_weightRead_7_data[1623 : 1616];
  assign dSP_1003_d = loadWeight_1_weightRead_7_data[1751 : 1744];
  assign dSP_1003_b = _zz_b_7[87 : 80];
  assign dSP_1004_a = loadWeight_1_weightRead_7_data[1631 : 1624];
  assign dSP_1004_d = loadWeight_1_weightRead_7_data[1759 : 1752];
  assign dSP_1004_b = _zz_b_7[95 : 88];
  assign dSP_1005_a = loadWeight_1_weightRead_7_data[1639 : 1632];
  assign dSP_1005_d = loadWeight_1_weightRead_7_data[1767 : 1760];
  assign dSP_1005_b = _zz_b_7[103 : 96];
  assign dSP_1006_a = loadWeight_1_weightRead_7_data[1647 : 1640];
  assign dSP_1006_d = loadWeight_1_weightRead_7_data[1775 : 1768];
  assign dSP_1006_b = _zz_b_7[111 : 104];
  assign dSP_1007_a = loadWeight_1_weightRead_7_data[1655 : 1648];
  assign dSP_1007_d = loadWeight_1_weightRead_7_data[1783 : 1776];
  assign dSP_1007_b = _zz_b_7[119 : 112];
  assign dSP_1008_a = loadWeight_1_weightRead_7_data[1663 : 1656];
  assign dSP_1008_d = loadWeight_1_weightRead_7_data[1791 : 1784];
  assign dSP_1008_b = _zz_b_7[127 : 120];
  assign dSP_1009_a = loadWeight_1_weightRead_7_data[1799 : 1792];
  assign dSP_1009_d = loadWeight_1_weightRead_7_data[1927 : 1920];
  assign dSP_1009_b = _zz_b_7[7 : 0];
  assign dSP_1010_a = loadWeight_1_weightRead_7_data[1807 : 1800];
  assign dSP_1010_d = loadWeight_1_weightRead_7_data[1935 : 1928];
  assign dSP_1010_b = _zz_b_7[15 : 8];
  assign dSP_1011_a = loadWeight_1_weightRead_7_data[1815 : 1808];
  assign dSP_1011_d = loadWeight_1_weightRead_7_data[1943 : 1936];
  assign dSP_1011_b = _zz_b_7[23 : 16];
  assign dSP_1012_a = loadWeight_1_weightRead_7_data[1823 : 1816];
  assign dSP_1012_d = loadWeight_1_weightRead_7_data[1951 : 1944];
  assign dSP_1012_b = _zz_b_7[31 : 24];
  assign dSP_1013_a = loadWeight_1_weightRead_7_data[1831 : 1824];
  assign dSP_1013_d = loadWeight_1_weightRead_7_data[1959 : 1952];
  assign dSP_1013_b = _zz_b_7[39 : 32];
  assign dSP_1014_a = loadWeight_1_weightRead_7_data[1839 : 1832];
  assign dSP_1014_d = loadWeight_1_weightRead_7_data[1967 : 1960];
  assign dSP_1014_b = _zz_b_7[47 : 40];
  assign dSP_1015_a = loadWeight_1_weightRead_7_data[1847 : 1840];
  assign dSP_1015_d = loadWeight_1_weightRead_7_data[1975 : 1968];
  assign dSP_1015_b = _zz_b_7[55 : 48];
  assign dSP_1016_a = loadWeight_1_weightRead_7_data[1855 : 1848];
  assign dSP_1016_d = loadWeight_1_weightRead_7_data[1983 : 1976];
  assign dSP_1016_b = _zz_b_7[63 : 56];
  assign dSP_1017_a = loadWeight_1_weightRead_7_data[1863 : 1856];
  assign dSP_1017_d = loadWeight_1_weightRead_7_data[1991 : 1984];
  assign dSP_1017_b = _zz_b_7[71 : 64];
  assign dSP_1018_a = loadWeight_1_weightRead_7_data[1871 : 1864];
  assign dSP_1018_d = loadWeight_1_weightRead_7_data[1999 : 1992];
  assign dSP_1018_b = _zz_b_7[79 : 72];
  assign dSP_1019_a = loadWeight_1_weightRead_7_data[1879 : 1872];
  assign dSP_1019_d = loadWeight_1_weightRead_7_data[2007 : 2000];
  assign dSP_1019_b = _zz_b_7[87 : 80];
  assign dSP_1020_a = loadWeight_1_weightRead_7_data[1887 : 1880];
  assign dSP_1020_d = loadWeight_1_weightRead_7_data[2015 : 2008];
  assign dSP_1020_b = _zz_b_7[95 : 88];
  assign dSP_1021_a = loadWeight_1_weightRead_7_data[1895 : 1888];
  assign dSP_1021_d = loadWeight_1_weightRead_7_data[2023 : 2016];
  assign dSP_1021_b = _zz_b_7[103 : 96];
  assign dSP_1022_a = loadWeight_1_weightRead_7_data[1903 : 1896];
  assign dSP_1022_d = loadWeight_1_weightRead_7_data[2031 : 2024];
  assign dSP_1022_b = _zz_b_7[111 : 104];
  assign dSP_1023_a = loadWeight_1_weightRead_7_data[1911 : 1904];
  assign dSP_1023_d = loadWeight_1_weightRead_7_data[2039 : 2032];
  assign dSP_1023_b = _zz_b_7[119 : 112];
  assign dSP_1024_a = loadWeight_1_weightRead_7_data[1919 : 1912];
  assign dSP_1024_d = loadWeight_1_weightRead_7_data[2047 : 2040];
  assign dSP_1024_b = _zz_b_7[127 : 120];
  assign dSP_1025_a = loadWeight_1_weightRead_8_data[7 : 0];
  assign dSP_1025_d = loadWeight_1_weightRead_8_data[135 : 128];
  assign dSP_1025_b = _zz_b_8[7 : 0];
  assign dSP_1026_a = loadWeight_1_weightRead_8_data[15 : 8];
  assign dSP_1026_d = loadWeight_1_weightRead_8_data[143 : 136];
  assign dSP_1026_b = _zz_b_8[15 : 8];
  assign dSP_1027_a = loadWeight_1_weightRead_8_data[23 : 16];
  assign dSP_1027_d = loadWeight_1_weightRead_8_data[151 : 144];
  assign dSP_1027_b = _zz_b_8[23 : 16];
  assign dSP_1028_a = loadWeight_1_weightRead_8_data[31 : 24];
  assign dSP_1028_d = loadWeight_1_weightRead_8_data[159 : 152];
  assign dSP_1028_b = _zz_b_8[31 : 24];
  assign dSP_1029_a = loadWeight_1_weightRead_8_data[39 : 32];
  assign dSP_1029_d = loadWeight_1_weightRead_8_data[167 : 160];
  assign dSP_1029_b = _zz_b_8[39 : 32];
  assign dSP_1030_a = loadWeight_1_weightRead_8_data[47 : 40];
  assign dSP_1030_d = loadWeight_1_weightRead_8_data[175 : 168];
  assign dSP_1030_b = _zz_b_8[47 : 40];
  assign dSP_1031_a = loadWeight_1_weightRead_8_data[55 : 48];
  assign dSP_1031_d = loadWeight_1_weightRead_8_data[183 : 176];
  assign dSP_1031_b = _zz_b_8[55 : 48];
  assign dSP_1032_a = loadWeight_1_weightRead_8_data[63 : 56];
  assign dSP_1032_d = loadWeight_1_weightRead_8_data[191 : 184];
  assign dSP_1032_b = _zz_b_8[63 : 56];
  assign dSP_1033_a = loadWeight_1_weightRead_8_data[71 : 64];
  assign dSP_1033_d = loadWeight_1_weightRead_8_data[199 : 192];
  assign dSP_1033_b = _zz_b_8[71 : 64];
  assign dSP_1034_a = loadWeight_1_weightRead_8_data[79 : 72];
  assign dSP_1034_d = loadWeight_1_weightRead_8_data[207 : 200];
  assign dSP_1034_b = _zz_b_8[79 : 72];
  assign dSP_1035_a = loadWeight_1_weightRead_8_data[87 : 80];
  assign dSP_1035_d = loadWeight_1_weightRead_8_data[215 : 208];
  assign dSP_1035_b = _zz_b_8[87 : 80];
  assign dSP_1036_a = loadWeight_1_weightRead_8_data[95 : 88];
  assign dSP_1036_d = loadWeight_1_weightRead_8_data[223 : 216];
  assign dSP_1036_b = _zz_b_8[95 : 88];
  assign dSP_1037_a = loadWeight_1_weightRead_8_data[103 : 96];
  assign dSP_1037_d = loadWeight_1_weightRead_8_data[231 : 224];
  assign dSP_1037_b = _zz_b_8[103 : 96];
  assign dSP_1038_a = loadWeight_1_weightRead_8_data[111 : 104];
  assign dSP_1038_d = loadWeight_1_weightRead_8_data[239 : 232];
  assign dSP_1038_b = _zz_b_8[111 : 104];
  assign dSP_1039_a = loadWeight_1_weightRead_8_data[119 : 112];
  assign dSP_1039_d = loadWeight_1_weightRead_8_data[247 : 240];
  assign dSP_1039_b = _zz_b_8[119 : 112];
  assign dSP_1040_a = loadWeight_1_weightRead_8_data[127 : 120];
  assign dSP_1040_d = loadWeight_1_weightRead_8_data[255 : 248];
  assign dSP_1040_b = _zz_b_8[127 : 120];
  assign dSP_1041_a = loadWeight_1_weightRead_8_data[263 : 256];
  assign dSP_1041_d = loadWeight_1_weightRead_8_data[391 : 384];
  assign dSP_1041_b = _zz_b_8[7 : 0];
  assign dSP_1042_a = loadWeight_1_weightRead_8_data[271 : 264];
  assign dSP_1042_d = loadWeight_1_weightRead_8_data[399 : 392];
  assign dSP_1042_b = _zz_b_8[15 : 8];
  assign dSP_1043_a = loadWeight_1_weightRead_8_data[279 : 272];
  assign dSP_1043_d = loadWeight_1_weightRead_8_data[407 : 400];
  assign dSP_1043_b = _zz_b_8[23 : 16];
  assign dSP_1044_a = loadWeight_1_weightRead_8_data[287 : 280];
  assign dSP_1044_d = loadWeight_1_weightRead_8_data[415 : 408];
  assign dSP_1044_b = _zz_b_8[31 : 24];
  assign dSP_1045_a = loadWeight_1_weightRead_8_data[295 : 288];
  assign dSP_1045_d = loadWeight_1_weightRead_8_data[423 : 416];
  assign dSP_1045_b = _zz_b_8[39 : 32];
  assign dSP_1046_a = loadWeight_1_weightRead_8_data[303 : 296];
  assign dSP_1046_d = loadWeight_1_weightRead_8_data[431 : 424];
  assign dSP_1046_b = _zz_b_8[47 : 40];
  assign dSP_1047_a = loadWeight_1_weightRead_8_data[311 : 304];
  assign dSP_1047_d = loadWeight_1_weightRead_8_data[439 : 432];
  assign dSP_1047_b = _zz_b_8[55 : 48];
  assign dSP_1048_a = loadWeight_1_weightRead_8_data[319 : 312];
  assign dSP_1048_d = loadWeight_1_weightRead_8_data[447 : 440];
  assign dSP_1048_b = _zz_b_8[63 : 56];
  assign dSP_1049_a = loadWeight_1_weightRead_8_data[327 : 320];
  assign dSP_1049_d = loadWeight_1_weightRead_8_data[455 : 448];
  assign dSP_1049_b = _zz_b_8[71 : 64];
  assign dSP_1050_a = loadWeight_1_weightRead_8_data[335 : 328];
  assign dSP_1050_d = loadWeight_1_weightRead_8_data[463 : 456];
  assign dSP_1050_b = _zz_b_8[79 : 72];
  assign dSP_1051_a = loadWeight_1_weightRead_8_data[343 : 336];
  assign dSP_1051_d = loadWeight_1_weightRead_8_data[471 : 464];
  assign dSP_1051_b = _zz_b_8[87 : 80];
  assign dSP_1052_a = loadWeight_1_weightRead_8_data[351 : 344];
  assign dSP_1052_d = loadWeight_1_weightRead_8_data[479 : 472];
  assign dSP_1052_b = _zz_b_8[95 : 88];
  assign dSP_1053_a = loadWeight_1_weightRead_8_data[359 : 352];
  assign dSP_1053_d = loadWeight_1_weightRead_8_data[487 : 480];
  assign dSP_1053_b = _zz_b_8[103 : 96];
  assign dSP_1054_a = loadWeight_1_weightRead_8_data[367 : 360];
  assign dSP_1054_d = loadWeight_1_weightRead_8_data[495 : 488];
  assign dSP_1054_b = _zz_b_8[111 : 104];
  assign dSP_1055_a = loadWeight_1_weightRead_8_data[375 : 368];
  assign dSP_1055_d = loadWeight_1_weightRead_8_data[503 : 496];
  assign dSP_1055_b = _zz_b_8[119 : 112];
  assign dSP_1056_a = loadWeight_1_weightRead_8_data[383 : 376];
  assign dSP_1056_d = loadWeight_1_weightRead_8_data[511 : 504];
  assign dSP_1056_b = _zz_b_8[127 : 120];
  assign dSP_1057_a = loadWeight_1_weightRead_8_data[519 : 512];
  assign dSP_1057_d = loadWeight_1_weightRead_8_data[647 : 640];
  assign dSP_1057_b = _zz_b_8[7 : 0];
  assign dSP_1058_a = loadWeight_1_weightRead_8_data[527 : 520];
  assign dSP_1058_d = loadWeight_1_weightRead_8_data[655 : 648];
  assign dSP_1058_b = _zz_b_8[15 : 8];
  assign dSP_1059_a = loadWeight_1_weightRead_8_data[535 : 528];
  assign dSP_1059_d = loadWeight_1_weightRead_8_data[663 : 656];
  assign dSP_1059_b = _zz_b_8[23 : 16];
  assign dSP_1060_a = loadWeight_1_weightRead_8_data[543 : 536];
  assign dSP_1060_d = loadWeight_1_weightRead_8_data[671 : 664];
  assign dSP_1060_b = _zz_b_8[31 : 24];
  assign dSP_1061_a = loadWeight_1_weightRead_8_data[551 : 544];
  assign dSP_1061_d = loadWeight_1_weightRead_8_data[679 : 672];
  assign dSP_1061_b = _zz_b_8[39 : 32];
  assign dSP_1062_a = loadWeight_1_weightRead_8_data[559 : 552];
  assign dSP_1062_d = loadWeight_1_weightRead_8_data[687 : 680];
  assign dSP_1062_b = _zz_b_8[47 : 40];
  assign dSP_1063_a = loadWeight_1_weightRead_8_data[567 : 560];
  assign dSP_1063_d = loadWeight_1_weightRead_8_data[695 : 688];
  assign dSP_1063_b = _zz_b_8[55 : 48];
  assign dSP_1064_a = loadWeight_1_weightRead_8_data[575 : 568];
  assign dSP_1064_d = loadWeight_1_weightRead_8_data[703 : 696];
  assign dSP_1064_b = _zz_b_8[63 : 56];
  assign dSP_1065_a = loadWeight_1_weightRead_8_data[583 : 576];
  assign dSP_1065_d = loadWeight_1_weightRead_8_data[711 : 704];
  assign dSP_1065_b = _zz_b_8[71 : 64];
  assign dSP_1066_a = loadWeight_1_weightRead_8_data[591 : 584];
  assign dSP_1066_d = loadWeight_1_weightRead_8_data[719 : 712];
  assign dSP_1066_b = _zz_b_8[79 : 72];
  assign dSP_1067_a = loadWeight_1_weightRead_8_data[599 : 592];
  assign dSP_1067_d = loadWeight_1_weightRead_8_data[727 : 720];
  assign dSP_1067_b = _zz_b_8[87 : 80];
  assign dSP_1068_a = loadWeight_1_weightRead_8_data[607 : 600];
  assign dSP_1068_d = loadWeight_1_weightRead_8_data[735 : 728];
  assign dSP_1068_b = _zz_b_8[95 : 88];
  assign dSP_1069_a = loadWeight_1_weightRead_8_data[615 : 608];
  assign dSP_1069_d = loadWeight_1_weightRead_8_data[743 : 736];
  assign dSP_1069_b = _zz_b_8[103 : 96];
  assign dSP_1070_a = loadWeight_1_weightRead_8_data[623 : 616];
  assign dSP_1070_d = loadWeight_1_weightRead_8_data[751 : 744];
  assign dSP_1070_b = _zz_b_8[111 : 104];
  assign dSP_1071_a = loadWeight_1_weightRead_8_data[631 : 624];
  assign dSP_1071_d = loadWeight_1_weightRead_8_data[759 : 752];
  assign dSP_1071_b = _zz_b_8[119 : 112];
  assign dSP_1072_a = loadWeight_1_weightRead_8_data[639 : 632];
  assign dSP_1072_d = loadWeight_1_weightRead_8_data[767 : 760];
  assign dSP_1072_b = _zz_b_8[127 : 120];
  assign dSP_1073_a = loadWeight_1_weightRead_8_data[775 : 768];
  assign dSP_1073_d = loadWeight_1_weightRead_8_data[903 : 896];
  assign dSP_1073_b = _zz_b_8[7 : 0];
  assign dSP_1074_a = loadWeight_1_weightRead_8_data[783 : 776];
  assign dSP_1074_d = loadWeight_1_weightRead_8_data[911 : 904];
  assign dSP_1074_b = _zz_b_8[15 : 8];
  assign dSP_1075_a = loadWeight_1_weightRead_8_data[791 : 784];
  assign dSP_1075_d = loadWeight_1_weightRead_8_data[919 : 912];
  assign dSP_1075_b = _zz_b_8[23 : 16];
  assign dSP_1076_a = loadWeight_1_weightRead_8_data[799 : 792];
  assign dSP_1076_d = loadWeight_1_weightRead_8_data[927 : 920];
  assign dSP_1076_b = _zz_b_8[31 : 24];
  assign dSP_1077_a = loadWeight_1_weightRead_8_data[807 : 800];
  assign dSP_1077_d = loadWeight_1_weightRead_8_data[935 : 928];
  assign dSP_1077_b = _zz_b_8[39 : 32];
  assign dSP_1078_a = loadWeight_1_weightRead_8_data[815 : 808];
  assign dSP_1078_d = loadWeight_1_weightRead_8_data[943 : 936];
  assign dSP_1078_b = _zz_b_8[47 : 40];
  assign dSP_1079_a = loadWeight_1_weightRead_8_data[823 : 816];
  assign dSP_1079_d = loadWeight_1_weightRead_8_data[951 : 944];
  assign dSP_1079_b = _zz_b_8[55 : 48];
  assign dSP_1080_a = loadWeight_1_weightRead_8_data[831 : 824];
  assign dSP_1080_d = loadWeight_1_weightRead_8_data[959 : 952];
  assign dSP_1080_b = _zz_b_8[63 : 56];
  assign dSP_1081_a = loadWeight_1_weightRead_8_data[839 : 832];
  assign dSP_1081_d = loadWeight_1_weightRead_8_data[967 : 960];
  assign dSP_1081_b = _zz_b_8[71 : 64];
  assign dSP_1082_a = loadWeight_1_weightRead_8_data[847 : 840];
  assign dSP_1082_d = loadWeight_1_weightRead_8_data[975 : 968];
  assign dSP_1082_b = _zz_b_8[79 : 72];
  assign dSP_1083_a = loadWeight_1_weightRead_8_data[855 : 848];
  assign dSP_1083_d = loadWeight_1_weightRead_8_data[983 : 976];
  assign dSP_1083_b = _zz_b_8[87 : 80];
  assign dSP_1084_a = loadWeight_1_weightRead_8_data[863 : 856];
  assign dSP_1084_d = loadWeight_1_weightRead_8_data[991 : 984];
  assign dSP_1084_b = _zz_b_8[95 : 88];
  assign dSP_1085_a = loadWeight_1_weightRead_8_data[871 : 864];
  assign dSP_1085_d = loadWeight_1_weightRead_8_data[999 : 992];
  assign dSP_1085_b = _zz_b_8[103 : 96];
  assign dSP_1086_a = loadWeight_1_weightRead_8_data[879 : 872];
  assign dSP_1086_d = loadWeight_1_weightRead_8_data[1007 : 1000];
  assign dSP_1086_b = _zz_b_8[111 : 104];
  assign dSP_1087_a = loadWeight_1_weightRead_8_data[887 : 880];
  assign dSP_1087_d = loadWeight_1_weightRead_8_data[1015 : 1008];
  assign dSP_1087_b = _zz_b_8[119 : 112];
  assign dSP_1088_a = loadWeight_1_weightRead_8_data[895 : 888];
  assign dSP_1088_d = loadWeight_1_weightRead_8_data[1023 : 1016];
  assign dSP_1088_b = _zz_b_8[127 : 120];
  assign dSP_1089_a = loadWeight_1_weightRead_8_data[1031 : 1024];
  assign dSP_1089_d = loadWeight_1_weightRead_8_data[1159 : 1152];
  assign dSP_1089_b = _zz_b_8[7 : 0];
  assign dSP_1090_a = loadWeight_1_weightRead_8_data[1039 : 1032];
  assign dSP_1090_d = loadWeight_1_weightRead_8_data[1167 : 1160];
  assign dSP_1090_b = _zz_b_8[15 : 8];
  assign dSP_1091_a = loadWeight_1_weightRead_8_data[1047 : 1040];
  assign dSP_1091_d = loadWeight_1_weightRead_8_data[1175 : 1168];
  assign dSP_1091_b = _zz_b_8[23 : 16];
  assign dSP_1092_a = loadWeight_1_weightRead_8_data[1055 : 1048];
  assign dSP_1092_d = loadWeight_1_weightRead_8_data[1183 : 1176];
  assign dSP_1092_b = _zz_b_8[31 : 24];
  assign dSP_1093_a = loadWeight_1_weightRead_8_data[1063 : 1056];
  assign dSP_1093_d = loadWeight_1_weightRead_8_data[1191 : 1184];
  assign dSP_1093_b = _zz_b_8[39 : 32];
  assign dSP_1094_a = loadWeight_1_weightRead_8_data[1071 : 1064];
  assign dSP_1094_d = loadWeight_1_weightRead_8_data[1199 : 1192];
  assign dSP_1094_b = _zz_b_8[47 : 40];
  assign dSP_1095_a = loadWeight_1_weightRead_8_data[1079 : 1072];
  assign dSP_1095_d = loadWeight_1_weightRead_8_data[1207 : 1200];
  assign dSP_1095_b = _zz_b_8[55 : 48];
  assign dSP_1096_a = loadWeight_1_weightRead_8_data[1087 : 1080];
  assign dSP_1096_d = loadWeight_1_weightRead_8_data[1215 : 1208];
  assign dSP_1096_b = _zz_b_8[63 : 56];
  assign dSP_1097_a = loadWeight_1_weightRead_8_data[1095 : 1088];
  assign dSP_1097_d = loadWeight_1_weightRead_8_data[1223 : 1216];
  assign dSP_1097_b = _zz_b_8[71 : 64];
  assign dSP_1098_a = loadWeight_1_weightRead_8_data[1103 : 1096];
  assign dSP_1098_d = loadWeight_1_weightRead_8_data[1231 : 1224];
  assign dSP_1098_b = _zz_b_8[79 : 72];
  assign dSP_1099_a = loadWeight_1_weightRead_8_data[1111 : 1104];
  assign dSP_1099_d = loadWeight_1_weightRead_8_data[1239 : 1232];
  assign dSP_1099_b = _zz_b_8[87 : 80];
  assign dSP_1100_a = loadWeight_1_weightRead_8_data[1119 : 1112];
  assign dSP_1100_d = loadWeight_1_weightRead_8_data[1247 : 1240];
  assign dSP_1100_b = _zz_b_8[95 : 88];
  assign dSP_1101_a = loadWeight_1_weightRead_8_data[1127 : 1120];
  assign dSP_1101_d = loadWeight_1_weightRead_8_data[1255 : 1248];
  assign dSP_1101_b = _zz_b_8[103 : 96];
  assign dSP_1102_a = loadWeight_1_weightRead_8_data[1135 : 1128];
  assign dSP_1102_d = loadWeight_1_weightRead_8_data[1263 : 1256];
  assign dSP_1102_b = _zz_b_8[111 : 104];
  assign dSP_1103_a = loadWeight_1_weightRead_8_data[1143 : 1136];
  assign dSP_1103_d = loadWeight_1_weightRead_8_data[1271 : 1264];
  assign dSP_1103_b = _zz_b_8[119 : 112];
  assign dSP_1104_a = loadWeight_1_weightRead_8_data[1151 : 1144];
  assign dSP_1104_d = loadWeight_1_weightRead_8_data[1279 : 1272];
  assign dSP_1104_b = _zz_b_8[127 : 120];
  assign dSP_1105_a = loadWeight_1_weightRead_8_data[1287 : 1280];
  assign dSP_1105_d = loadWeight_1_weightRead_8_data[1415 : 1408];
  assign dSP_1105_b = _zz_b_8[7 : 0];
  assign dSP_1106_a = loadWeight_1_weightRead_8_data[1295 : 1288];
  assign dSP_1106_d = loadWeight_1_weightRead_8_data[1423 : 1416];
  assign dSP_1106_b = _zz_b_8[15 : 8];
  assign dSP_1107_a = loadWeight_1_weightRead_8_data[1303 : 1296];
  assign dSP_1107_d = loadWeight_1_weightRead_8_data[1431 : 1424];
  assign dSP_1107_b = _zz_b_8[23 : 16];
  assign dSP_1108_a = loadWeight_1_weightRead_8_data[1311 : 1304];
  assign dSP_1108_d = loadWeight_1_weightRead_8_data[1439 : 1432];
  assign dSP_1108_b = _zz_b_8[31 : 24];
  assign dSP_1109_a = loadWeight_1_weightRead_8_data[1319 : 1312];
  assign dSP_1109_d = loadWeight_1_weightRead_8_data[1447 : 1440];
  assign dSP_1109_b = _zz_b_8[39 : 32];
  assign dSP_1110_a = loadWeight_1_weightRead_8_data[1327 : 1320];
  assign dSP_1110_d = loadWeight_1_weightRead_8_data[1455 : 1448];
  assign dSP_1110_b = _zz_b_8[47 : 40];
  assign dSP_1111_a = loadWeight_1_weightRead_8_data[1335 : 1328];
  assign dSP_1111_d = loadWeight_1_weightRead_8_data[1463 : 1456];
  assign dSP_1111_b = _zz_b_8[55 : 48];
  assign dSP_1112_a = loadWeight_1_weightRead_8_data[1343 : 1336];
  assign dSP_1112_d = loadWeight_1_weightRead_8_data[1471 : 1464];
  assign dSP_1112_b = _zz_b_8[63 : 56];
  assign dSP_1113_a = loadWeight_1_weightRead_8_data[1351 : 1344];
  assign dSP_1113_d = loadWeight_1_weightRead_8_data[1479 : 1472];
  assign dSP_1113_b = _zz_b_8[71 : 64];
  assign dSP_1114_a = loadWeight_1_weightRead_8_data[1359 : 1352];
  assign dSP_1114_d = loadWeight_1_weightRead_8_data[1487 : 1480];
  assign dSP_1114_b = _zz_b_8[79 : 72];
  assign dSP_1115_a = loadWeight_1_weightRead_8_data[1367 : 1360];
  assign dSP_1115_d = loadWeight_1_weightRead_8_data[1495 : 1488];
  assign dSP_1115_b = _zz_b_8[87 : 80];
  assign dSP_1116_a = loadWeight_1_weightRead_8_data[1375 : 1368];
  assign dSP_1116_d = loadWeight_1_weightRead_8_data[1503 : 1496];
  assign dSP_1116_b = _zz_b_8[95 : 88];
  assign dSP_1117_a = loadWeight_1_weightRead_8_data[1383 : 1376];
  assign dSP_1117_d = loadWeight_1_weightRead_8_data[1511 : 1504];
  assign dSP_1117_b = _zz_b_8[103 : 96];
  assign dSP_1118_a = loadWeight_1_weightRead_8_data[1391 : 1384];
  assign dSP_1118_d = loadWeight_1_weightRead_8_data[1519 : 1512];
  assign dSP_1118_b = _zz_b_8[111 : 104];
  assign dSP_1119_a = loadWeight_1_weightRead_8_data[1399 : 1392];
  assign dSP_1119_d = loadWeight_1_weightRead_8_data[1527 : 1520];
  assign dSP_1119_b = _zz_b_8[119 : 112];
  assign dSP_1120_a = loadWeight_1_weightRead_8_data[1407 : 1400];
  assign dSP_1120_d = loadWeight_1_weightRead_8_data[1535 : 1528];
  assign dSP_1120_b = _zz_b_8[127 : 120];
  assign dSP_1121_a = loadWeight_1_weightRead_8_data[1543 : 1536];
  assign dSP_1121_d = loadWeight_1_weightRead_8_data[1671 : 1664];
  assign dSP_1121_b = _zz_b_8[7 : 0];
  assign dSP_1122_a = loadWeight_1_weightRead_8_data[1551 : 1544];
  assign dSP_1122_d = loadWeight_1_weightRead_8_data[1679 : 1672];
  assign dSP_1122_b = _zz_b_8[15 : 8];
  assign dSP_1123_a = loadWeight_1_weightRead_8_data[1559 : 1552];
  assign dSP_1123_d = loadWeight_1_weightRead_8_data[1687 : 1680];
  assign dSP_1123_b = _zz_b_8[23 : 16];
  assign dSP_1124_a = loadWeight_1_weightRead_8_data[1567 : 1560];
  assign dSP_1124_d = loadWeight_1_weightRead_8_data[1695 : 1688];
  assign dSP_1124_b = _zz_b_8[31 : 24];
  assign dSP_1125_a = loadWeight_1_weightRead_8_data[1575 : 1568];
  assign dSP_1125_d = loadWeight_1_weightRead_8_data[1703 : 1696];
  assign dSP_1125_b = _zz_b_8[39 : 32];
  assign dSP_1126_a = loadWeight_1_weightRead_8_data[1583 : 1576];
  assign dSP_1126_d = loadWeight_1_weightRead_8_data[1711 : 1704];
  assign dSP_1126_b = _zz_b_8[47 : 40];
  assign dSP_1127_a = loadWeight_1_weightRead_8_data[1591 : 1584];
  assign dSP_1127_d = loadWeight_1_weightRead_8_data[1719 : 1712];
  assign dSP_1127_b = _zz_b_8[55 : 48];
  assign dSP_1128_a = loadWeight_1_weightRead_8_data[1599 : 1592];
  assign dSP_1128_d = loadWeight_1_weightRead_8_data[1727 : 1720];
  assign dSP_1128_b = _zz_b_8[63 : 56];
  assign dSP_1129_a = loadWeight_1_weightRead_8_data[1607 : 1600];
  assign dSP_1129_d = loadWeight_1_weightRead_8_data[1735 : 1728];
  assign dSP_1129_b = _zz_b_8[71 : 64];
  assign dSP_1130_a = loadWeight_1_weightRead_8_data[1615 : 1608];
  assign dSP_1130_d = loadWeight_1_weightRead_8_data[1743 : 1736];
  assign dSP_1130_b = _zz_b_8[79 : 72];
  assign dSP_1131_a = loadWeight_1_weightRead_8_data[1623 : 1616];
  assign dSP_1131_d = loadWeight_1_weightRead_8_data[1751 : 1744];
  assign dSP_1131_b = _zz_b_8[87 : 80];
  assign dSP_1132_a = loadWeight_1_weightRead_8_data[1631 : 1624];
  assign dSP_1132_d = loadWeight_1_weightRead_8_data[1759 : 1752];
  assign dSP_1132_b = _zz_b_8[95 : 88];
  assign dSP_1133_a = loadWeight_1_weightRead_8_data[1639 : 1632];
  assign dSP_1133_d = loadWeight_1_weightRead_8_data[1767 : 1760];
  assign dSP_1133_b = _zz_b_8[103 : 96];
  assign dSP_1134_a = loadWeight_1_weightRead_8_data[1647 : 1640];
  assign dSP_1134_d = loadWeight_1_weightRead_8_data[1775 : 1768];
  assign dSP_1134_b = _zz_b_8[111 : 104];
  assign dSP_1135_a = loadWeight_1_weightRead_8_data[1655 : 1648];
  assign dSP_1135_d = loadWeight_1_weightRead_8_data[1783 : 1776];
  assign dSP_1135_b = _zz_b_8[119 : 112];
  assign dSP_1136_a = loadWeight_1_weightRead_8_data[1663 : 1656];
  assign dSP_1136_d = loadWeight_1_weightRead_8_data[1791 : 1784];
  assign dSP_1136_b = _zz_b_8[127 : 120];
  assign dSP_1137_a = loadWeight_1_weightRead_8_data[1799 : 1792];
  assign dSP_1137_d = loadWeight_1_weightRead_8_data[1927 : 1920];
  assign dSP_1137_b = _zz_b_8[7 : 0];
  assign dSP_1138_a = loadWeight_1_weightRead_8_data[1807 : 1800];
  assign dSP_1138_d = loadWeight_1_weightRead_8_data[1935 : 1928];
  assign dSP_1138_b = _zz_b_8[15 : 8];
  assign dSP_1139_a = loadWeight_1_weightRead_8_data[1815 : 1808];
  assign dSP_1139_d = loadWeight_1_weightRead_8_data[1943 : 1936];
  assign dSP_1139_b = _zz_b_8[23 : 16];
  assign dSP_1140_a = loadWeight_1_weightRead_8_data[1823 : 1816];
  assign dSP_1140_d = loadWeight_1_weightRead_8_data[1951 : 1944];
  assign dSP_1140_b = _zz_b_8[31 : 24];
  assign dSP_1141_a = loadWeight_1_weightRead_8_data[1831 : 1824];
  assign dSP_1141_d = loadWeight_1_weightRead_8_data[1959 : 1952];
  assign dSP_1141_b = _zz_b_8[39 : 32];
  assign dSP_1142_a = loadWeight_1_weightRead_8_data[1839 : 1832];
  assign dSP_1142_d = loadWeight_1_weightRead_8_data[1967 : 1960];
  assign dSP_1142_b = _zz_b_8[47 : 40];
  assign dSP_1143_a = loadWeight_1_weightRead_8_data[1847 : 1840];
  assign dSP_1143_d = loadWeight_1_weightRead_8_data[1975 : 1968];
  assign dSP_1143_b = _zz_b_8[55 : 48];
  assign dSP_1144_a = loadWeight_1_weightRead_8_data[1855 : 1848];
  assign dSP_1144_d = loadWeight_1_weightRead_8_data[1983 : 1976];
  assign dSP_1144_b = _zz_b_8[63 : 56];
  assign dSP_1145_a = loadWeight_1_weightRead_8_data[1863 : 1856];
  assign dSP_1145_d = loadWeight_1_weightRead_8_data[1991 : 1984];
  assign dSP_1145_b = _zz_b_8[71 : 64];
  assign dSP_1146_a = loadWeight_1_weightRead_8_data[1871 : 1864];
  assign dSP_1146_d = loadWeight_1_weightRead_8_data[1999 : 1992];
  assign dSP_1146_b = _zz_b_8[79 : 72];
  assign dSP_1147_a = loadWeight_1_weightRead_8_data[1879 : 1872];
  assign dSP_1147_d = loadWeight_1_weightRead_8_data[2007 : 2000];
  assign dSP_1147_b = _zz_b_8[87 : 80];
  assign dSP_1148_a = loadWeight_1_weightRead_8_data[1887 : 1880];
  assign dSP_1148_d = loadWeight_1_weightRead_8_data[2015 : 2008];
  assign dSP_1148_b = _zz_b_8[95 : 88];
  assign dSP_1149_a = loadWeight_1_weightRead_8_data[1895 : 1888];
  assign dSP_1149_d = loadWeight_1_weightRead_8_data[2023 : 2016];
  assign dSP_1149_b = _zz_b_8[103 : 96];
  assign dSP_1150_a = loadWeight_1_weightRead_8_data[1903 : 1896];
  assign dSP_1150_d = loadWeight_1_weightRead_8_data[2031 : 2024];
  assign dSP_1150_b = _zz_b_8[111 : 104];
  assign dSP_1151_a = loadWeight_1_weightRead_8_data[1911 : 1904];
  assign dSP_1151_d = loadWeight_1_weightRead_8_data[2039 : 2032];
  assign dSP_1151_b = _zz_b_8[119 : 112];
  assign dSP_1152_a = loadWeight_1_weightRead_8_data[1919 : 1912];
  assign dSP_1152_d = loadWeight_1_weightRead_8_data[2047 : 2040];
  assign dSP_1152_b = _zz_b_8[127 : 120];
  assign addKernel_A_0 = dSP_1_p;
  assign addKernel_A_1 = dSP_129_p;
  assign addKernel_A_2 = dSP_257_p;
  assign addKernel_A_3 = dSP_385_p;
  assign addKernel_A_4 = dSP_513_p;
  assign addKernel_A_5 = dSP_641_p;
  assign addKernel_A_6 = dSP_769_p;
  assign addKernel_A_7 = dSP_897_p;
  assign addKernel_A_8 = dSP_1025_p;
  assign addKernel_1_A_0 = dSP_2_p;
  assign addKernel_1_A_1 = dSP_130_p;
  assign addKernel_1_A_2 = dSP_258_p;
  assign addKernel_1_A_3 = dSP_386_p;
  assign addKernel_1_A_4 = dSP_514_p;
  assign addKernel_1_A_5 = dSP_642_p;
  assign addKernel_1_A_6 = dSP_770_p;
  assign addKernel_1_A_7 = dSP_898_p;
  assign addKernel_1_A_8 = dSP_1026_p;
  assign addKernel_2_A_0 = dSP_3_p;
  assign addKernel_2_A_1 = dSP_131_p;
  assign addKernel_2_A_2 = dSP_259_p;
  assign addKernel_2_A_3 = dSP_387_p;
  assign addKernel_2_A_4 = dSP_515_p;
  assign addKernel_2_A_5 = dSP_643_p;
  assign addKernel_2_A_6 = dSP_771_p;
  assign addKernel_2_A_7 = dSP_899_p;
  assign addKernel_2_A_8 = dSP_1027_p;
  assign addKernel_3_A_0 = dSP_4_p;
  assign addKernel_3_A_1 = dSP_132_p;
  assign addKernel_3_A_2 = dSP_260_p;
  assign addKernel_3_A_3 = dSP_388_p;
  assign addKernel_3_A_4 = dSP_516_p;
  assign addKernel_3_A_5 = dSP_644_p;
  assign addKernel_3_A_6 = dSP_772_p;
  assign addKernel_3_A_7 = dSP_900_p;
  assign addKernel_3_A_8 = dSP_1028_p;
  assign addKernel_4_A_0 = dSP_5_p;
  assign addKernel_4_A_1 = dSP_133_p;
  assign addKernel_4_A_2 = dSP_261_p;
  assign addKernel_4_A_3 = dSP_389_p;
  assign addKernel_4_A_4 = dSP_517_p;
  assign addKernel_4_A_5 = dSP_645_p;
  assign addKernel_4_A_6 = dSP_773_p;
  assign addKernel_4_A_7 = dSP_901_p;
  assign addKernel_4_A_8 = dSP_1029_p;
  assign addKernel_5_A_0 = dSP_6_p;
  assign addKernel_5_A_1 = dSP_134_p;
  assign addKernel_5_A_2 = dSP_262_p;
  assign addKernel_5_A_3 = dSP_390_p;
  assign addKernel_5_A_4 = dSP_518_p;
  assign addKernel_5_A_5 = dSP_646_p;
  assign addKernel_5_A_6 = dSP_774_p;
  assign addKernel_5_A_7 = dSP_902_p;
  assign addKernel_5_A_8 = dSP_1030_p;
  assign addKernel_6_A_0 = dSP_7_p;
  assign addKernel_6_A_1 = dSP_135_p;
  assign addKernel_6_A_2 = dSP_263_p;
  assign addKernel_6_A_3 = dSP_391_p;
  assign addKernel_6_A_4 = dSP_519_p;
  assign addKernel_6_A_5 = dSP_647_p;
  assign addKernel_6_A_6 = dSP_775_p;
  assign addKernel_6_A_7 = dSP_903_p;
  assign addKernel_6_A_8 = dSP_1031_p;
  assign addKernel_7_A_0 = dSP_8_p;
  assign addKernel_7_A_1 = dSP_136_p;
  assign addKernel_7_A_2 = dSP_264_p;
  assign addKernel_7_A_3 = dSP_392_p;
  assign addKernel_7_A_4 = dSP_520_p;
  assign addKernel_7_A_5 = dSP_648_p;
  assign addKernel_7_A_6 = dSP_776_p;
  assign addKernel_7_A_7 = dSP_904_p;
  assign addKernel_7_A_8 = dSP_1032_p;
  assign addKernel_8_A_0 = dSP_9_p;
  assign addKernel_8_A_1 = dSP_137_p;
  assign addKernel_8_A_2 = dSP_265_p;
  assign addKernel_8_A_3 = dSP_393_p;
  assign addKernel_8_A_4 = dSP_521_p;
  assign addKernel_8_A_5 = dSP_649_p;
  assign addKernel_8_A_6 = dSP_777_p;
  assign addKernel_8_A_7 = dSP_905_p;
  assign addKernel_8_A_8 = dSP_1033_p;
  assign addKernel_9_A_0 = dSP_10_p;
  assign addKernel_9_A_1 = dSP_138_p;
  assign addKernel_9_A_2 = dSP_266_p;
  assign addKernel_9_A_3 = dSP_394_p;
  assign addKernel_9_A_4 = dSP_522_p;
  assign addKernel_9_A_5 = dSP_650_p;
  assign addKernel_9_A_6 = dSP_778_p;
  assign addKernel_9_A_7 = dSP_906_p;
  assign addKernel_9_A_8 = dSP_1034_p;
  assign addKernel_10_A_0 = dSP_11_p;
  assign addKernel_10_A_1 = dSP_139_p;
  assign addKernel_10_A_2 = dSP_267_p;
  assign addKernel_10_A_3 = dSP_395_p;
  assign addKernel_10_A_4 = dSP_523_p;
  assign addKernel_10_A_5 = dSP_651_p;
  assign addKernel_10_A_6 = dSP_779_p;
  assign addKernel_10_A_7 = dSP_907_p;
  assign addKernel_10_A_8 = dSP_1035_p;
  assign addKernel_11_A_0 = dSP_12_p;
  assign addKernel_11_A_1 = dSP_140_p;
  assign addKernel_11_A_2 = dSP_268_p;
  assign addKernel_11_A_3 = dSP_396_p;
  assign addKernel_11_A_4 = dSP_524_p;
  assign addKernel_11_A_5 = dSP_652_p;
  assign addKernel_11_A_6 = dSP_780_p;
  assign addKernel_11_A_7 = dSP_908_p;
  assign addKernel_11_A_8 = dSP_1036_p;
  assign addKernel_12_A_0 = dSP_13_p;
  assign addKernel_12_A_1 = dSP_141_p;
  assign addKernel_12_A_2 = dSP_269_p;
  assign addKernel_12_A_3 = dSP_397_p;
  assign addKernel_12_A_4 = dSP_525_p;
  assign addKernel_12_A_5 = dSP_653_p;
  assign addKernel_12_A_6 = dSP_781_p;
  assign addKernel_12_A_7 = dSP_909_p;
  assign addKernel_12_A_8 = dSP_1037_p;
  assign addKernel_13_A_0 = dSP_14_p;
  assign addKernel_13_A_1 = dSP_142_p;
  assign addKernel_13_A_2 = dSP_270_p;
  assign addKernel_13_A_3 = dSP_398_p;
  assign addKernel_13_A_4 = dSP_526_p;
  assign addKernel_13_A_5 = dSP_654_p;
  assign addKernel_13_A_6 = dSP_782_p;
  assign addKernel_13_A_7 = dSP_910_p;
  assign addKernel_13_A_8 = dSP_1038_p;
  assign addKernel_14_A_0 = dSP_15_p;
  assign addKernel_14_A_1 = dSP_143_p;
  assign addKernel_14_A_2 = dSP_271_p;
  assign addKernel_14_A_3 = dSP_399_p;
  assign addKernel_14_A_4 = dSP_527_p;
  assign addKernel_14_A_5 = dSP_655_p;
  assign addKernel_14_A_6 = dSP_783_p;
  assign addKernel_14_A_7 = dSP_911_p;
  assign addKernel_14_A_8 = dSP_1039_p;
  assign addKernel_15_A_0 = dSP_16_p;
  assign addKernel_15_A_1 = dSP_144_p;
  assign addKernel_15_A_2 = dSP_272_p;
  assign addKernel_15_A_3 = dSP_400_p;
  assign addKernel_15_A_4 = dSP_528_p;
  assign addKernel_15_A_5 = dSP_656_p;
  assign addKernel_15_A_6 = dSP_784_p;
  assign addKernel_15_A_7 = dSP_912_p;
  assign addKernel_15_A_8 = dSP_1040_p;
  assign addKernel_16_A_0 = dSP_17_p;
  assign addKernel_16_A_1 = dSP_145_p;
  assign addKernel_16_A_2 = dSP_273_p;
  assign addKernel_16_A_3 = dSP_401_p;
  assign addKernel_16_A_4 = dSP_529_p;
  assign addKernel_16_A_5 = dSP_657_p;
  assign addKernel_16_A_6 = dSP_785_p;
  assign addKernel_16_A_7 = dSP_913_p;
  assign addKernel_16_A_8 = dSP_1041_p;
  assign addKernel_17_A_0 = dSP_18_p;
  assign addKernel_17_A_1 = dSP_146_p;
  assign addKernel_17_A_2 = dSP_274_p;
  assign addKernel_17_A_3 = dSP_402_p;
  assign addKernel_17_A_4 = dSP_530_p;
  assign addKernel_17_A_5 = dSP_658_p;
  assign addKernel_17_A_6 = dSP_786_p;
  assign addKernel_17_A_7 = dSP_914_p;
  assign addKernel_17_A_8 = dSP_1042_p;
  assign addKernel_18_A_0 = dSP_19_p;
  assign addKernel_18_A_1 = dSP_147_p;
  assign addKernel_18_A_2 = dSP_275_p;
  assign addKernel_18_A_3 = dSP_403_p;
  assign addKernel_18_A_4 = dSP_531_p;
  assign addKernel_18_A_5 = dSP_659_p;
  assign addKernel_18_A_6 = dSP_787_p;
  assign addKernel_18_A_7 = dSP_915_p;
  assign addKernel_18_A_8 = dSP_1043_p;
  assign addKernel_19_A_0 = dSP_20_p;
  assign addKernel_19_A_1 = dSP_148_p;
  assign addKernel_19_A_2 = dSP_276_p;
  assign addKernel_19_A_3 = dSP_404_p;
  assign addKernel_19_A_4 = dSP_532_p;
  assign addKernel_19_A_5 = dSP_660_p;
  assign addKernel_19_A_6 = dSP_788_p;
  assign addKernel_19_A_7 = dSP_916_p;
  assign addKernel_19_A_8 = dSP_1044_p;
  assign addKernel_20_A_0 = dSP_21_p;
  assign addKernel_20_A_1 = dSP_149_p;
  assign addKernel_20_A_2 = dSP_277_p;
  assign addKernel_20_A_3 = dSP_405_p;
  assign addKernel_20_A_4 = dSP_533_p;
  assign addKernel_20_A_5 = dSP_661_p;
  assign addKernel_20_A_6 = dSP_789_p;
  assign addKernel_20_A_7 = dSP_917_p;
  assign addKernel_20_A_8 = dSP_1045_p;
  assign addKernel_21_A_0 = dSP_22_p;
  assign addKernel_21_A_1 = dSP_150_p;
  assign addKernel_21_A_2 = dSP_278_p;
  assign addKernel_21_A_3 = dSP_406_p;
  assign addKernel_21_A_4 = dSP_534_p;
  assign addKernel_21_A_5 = dSP_662_p;
  assign addKernel_21_A_6 = dSP_790_p;
  assign addKernel_21_A_7 = dSP_918_p;
  assign addKernel_21_A_8 = dSP_1046_p;
  assign addKernel_22_A_0 = dSP_23_p;
  assign addKernel_22_A_1 = dSP_151_p;
  assign addKernel_22_A_2 = dSP_279_p;
  assign addKernel_22_A_3 = dSP_407_p;
  assign addKernel_22_A_4 = dSP_535_p;
  assign addKernel_22_A_5 = dSP_663_p;
  assign addKernel_22_A_6 = dSP_791_p;
  assign addKernel_22_A_7 = dSP_919_p;
  assign addKernel_22_A_8 = dSP_1047_p;
  assign addKernel_23_A_0 = dSP_24_p;
  assign addKernel_23_A_1 = dSP_152_p;
  assign addKernel_23_A_2 = dSP_280_p;
  assign addKernel_23_A_3 = dSP_408_p;
  assign addKernel_23_A_4 = dSP_536_p;
  assign addKernel_23_A_5 = dSP_664_p;
  assign addKernel_23_A_6 = dSP_792_p;
  assign addKernel_23_A_7 = dSP_920_p;
  assign addKernel_23_A_8 = dSP_1048_p;
  assign addKernel_24_A_0 = dSP_25_p;
  assign addKernel_24_A_1 = dSP_153_p;
  assign addKernel_24_A_2 = dSP_281_p;
  assign addKernel_24_A_3 = dSP_409_p;
  assign addKernel_24_A_4 = dSP_537_p;
  assign addKernel_24_A_5 = dSP_665_p;
  assign addKernel_24_A_6 = dSP_793_p;
  assign addKernel_24_A_7 = dSP_921_p;
  assign addKernel_24_A_8 = dSP_1049_p;
  assign addKernel_25_A_0 = dSP_26_p;
  assign addKernel_25_A_1 = dSP_154_p;
  assign addKernel_25_A_2 = dSP_282_p;
  assign addKernel_25_A_3 = dSP_410_p;
  assign addKernel_25_A_4 = dSP_538_p;
  assign addKernel_25_A_5 = dSP_666_p;
  assign addKernel_25_A_6 = dSP_794_p;
  assign addKernel_25_A_7 = dSP_922_p;
  assign addKernel_25_A_8 = dSP_1050_p;
  assign addKernel_26_A_0 = dSP_27_p;
  assign addKernel_26_A_1 = dSP_155_p;
  assign addKernel_26_A_2 = dSP_283_p;
  assign addKernel_26_A_3 = dSP_411_p;
  assign addKernel_26_A_4 = dSP_539_p;
  assign addKernel_26_A_5 = dSP_667_p;
  assign addKernel_26_A_6 = dSP_795_p;
  assign addKernel_26_A_7 = dSP_923_p;
  assign addKernel_26_A_8 = dSP_1051_p;
  assign addKernel_27_A_0 = dSP_28_p;
  assign addKernel_27_A_1 = dSP_156_p;
  assign addKernel_27_A_2 = dSP_284_p;
  assign addKernel_27_A_3 = dSP_412_p;
  assign addKernel_27_A_4 = dSP_540_p;
  assign addKernel_27_A_5 = dSP_668_p;
  assign addKernel_27_A_6 = dSP_796_p;
  assign addKernel_27_A_7 = dSP_924_p;
  assign addKernel_27_A_8 = dSP_1052_p;
  assign addKernel_28_A_0 = dSP_29_p;
  assign addKernel_28_A_1 = dSP_157_p;
  assign addKernel_28_A_2 = dSP_285_p;
  assign addKernel_28_A_3 = dSP_413_p;
  assign addKernel_28_A_4 = dSP_541_p;
  assign addKernel_28_A_5 = dSP_669_p;
  assign addKernel_28_A_6 = dSP_797_p;
  assign addKernel_28_A_7 = dSP_925_p;
  assign addKernel_28_A_8 = dSP_1053_p;
  assign addKernel_29_A_0 = dSP_30_p;
  assign addKernel_29_A_1 = dSP_158_p;
  assign addKernel_29_A_2 = dSP_286_p;
  assign addKernel_29_A_3 = dSP_414_p;
  assign addKernel_29_A_4 = dSP_542_p;
  assign addKernel_29_A_5 = dSP_670_p;
  assign addKernel_29_A_6 = dSP_798_p;
  assign addKernel_29_A_7 = dSP_926_p;
  assign addKernel_29_A_8 = dSP_1054_p;
  assign addKernel_30_A_0 = dSP_31_p;
  assign addKernel_30_A_1 = dSP_159_p;
  assign addKernel_30_A_2 = dSP_287_p;
  assign addKernel_30_A_3 = dSP_415_p;
  assign addKernel_30_A_4 = dSP_543_p;
  assign addKernel_30_A_5 = dSP_671_p;
  assign addKernel_30_A_6 = dSP_799_p;
  assign addKernel_30_A_7 = dSP_927_p;
  assign addKernel_30_A_8 = dSP_1055_p;
  assign addKernel_31_A_0 = dSP_32_p;
  assign addKernel_31_A_1 = dSP_160_p;
  assign addKernel_31_A_2 = dSP_288_p;
  assign addKernel_31_A_3 = dSP_416_p;
  assign addKernel_31_A_4 = dSP_544_p;
  assign addKernel_31_A_5 = dSP_672_p;
  assign addKernel_31_A_6 = dSP_800_p;
  assign addKernel_31_A_7 = dSP_928_p;
  assign addKernel_31_A_8 = dSP_1056_p;
  assign addKernel_32_A_0 = dSP_33_p;
  assign addKernel_32_A_1 = dSP_161_p;
  assign addKernel_32_A_2 = dSP_289_p;
  assign addKernel_32_A_3 = dSP_417_p;
  assign addKernel_32_A_4 = dSP_545_p;
  assign addKernel_32_A_5 = dSP_673_p;
  assign addKernel_32_A_6 = dSP_801_p;
  assign addKernel_32_A_7 = dSP_929_p;
  assign addKernel_32_A_8 = dSP_1057_p;
  assign addKernel_33_A_0 = dSP_34_p;
  assign addKernel_33_A_1 = dSP_162_p;
  assign addKernel_33_A_2 = dSP_290_p;
  assign addKernel_33_A_3 = dSP_418_p;
  assign addKernel_33_A_4 = dSP_546_p;
  assign addKernel_33_A_5 = dSP_674_p;
  assign addKernel_33_A_6 = dSP_802_p;
  assign addKernel_33_A_7 = dSP_930_p;
  assign addKernel_33_A_8 = dSP_1058_p;
  assign addKernel_34_A_0 = dSP_35_p;
  assign addKernel_34_A_1 = dSP_163_p;
  assign addKernel_34_A_2 = dSP_291_p;
  assign addKernel_34_A_3 = dSP_419_p;
  assign addKernel_34_A_4 = dSP_547_p;
  assign addKernel_34_A_5 = dSP_675_p;
  assign addKernel_34_A_6 = dSP_803_p;
  assign addKernel_34_A_7 = dSP_931_p;
  assign addKernel_34_A_8 = dSP_1059_p;
  assign addKernel_35_A_0 = dSP_36_p;
  assign addKernel_35_A_1 = dSP_164_p;
  assign addKernel_35_A_2 = dSP_292_p;
  assign addKernel_35_A_3 = dSP_420_p;
  assign addKernel_35_A_4 = dSP_548_p;
  assign addKernel_35_A_5 = dSP_676_p;
  assign addKernel_35_A_6 = dSP_804_p;
  assign addKernel_35_A_7 = dSP_932_p;
  assign addKernel_35_A_8 = dSP_1060_p;
  assign addKernel_36_A_0 = dSP_37_p;
  assign addKernel_36_A_1 = dSP_165_p;
  assign addKernel_36_A_2 = dSP_293_p;
  assign addKernel_36_A_3 = dSP_421_p;
  assign addKernel_36_A_4 = dSP_549_p;
  assign addKernel_36_A_5 = dSP_677_p;
  assign addKernel_36_A_6 = dSP_805_p;
  assign addKernel_36_A_7 = dSP_933_p;
  assign addKernel_36_A_8 = dSP_1061_p;
  assign addKernel_37_A_0 = dSP_38_p;
  assign addKernel_37_A_1 = dSP_166_p;
  assign addKernel_37_A_2 = dSP_294_p;
  assign addKernel_37_A_3 = dSP_422_p;
  assign addKernel_37_A_4 = dSP_550_p;
  assign addKernel_37_A_5 = dSP_678_p;
  assign addKernel_37_A_6 = dSP_806_p;
  assign addKernel_37_A_7 = dSP_934_p;
  assign addKernel_37_A_8 = dSP_1062_p;
  assign addKernel_38_A_0 = dSP_39_p;
  assign addKernel_38_A_1 = dSP_167_p;
  assign addKernel_38_A_2 = dSP_295_p;
  assign addKernel_38_A_3 = dSP_423_p;
  assign addKernel_38_A_4 = dSP_551_p;
  assign addKernel_38_A_5 = dSP_679_p;
  assign addKernel_38_A_6 = dSP_807_p;
  assign addKernel_38_A_7 = dSP_935_p;
  assign addKernel_38_A_8 = dSP_1063_p;
  assign addKernel_39_A_0 = dSP_40_p;
  assign addKernel_39_A_1 = dSP_168_p;
  assign addKernel_39_A_2 = dSP_296_p;
  assign addKernel_39_A_3 = dSP_424_p;
  assign addKernel_39_A_4 = dSP_552_p;
  assign addKernel_39_A_5 = dSP_680_p;
  assign addKernel_39_A_6 = dSP_808_p;
  assign addKernel_39_A_7 = dSP_936_p;
  assign addKernel_39_A_8 = dSP_1064_p;
  assign addKernel_40_A_0 = dSP_41_p;
  assign addKernel_40_A_1 = dSP_169_p;
  assign addKernel_40_A_2 = dSP_297_p;
  assign addKernel_40_A_3 = dSP_425_p;
  assign addKernel_40_A_4 = dSP_553_p;
  assign addKernel_40_A_5 = dSP_681_p;
  assign addKernel_40_A_6 = dSP_809_p;
  assign addKernel_40_A_7 = dSP_937_p;
  assign addKernel_40_A_8 = dSP_1065_p;
  assign addKernel_41_A_0 = dSP_42_p;
  assign addKernel_41_A_1 = dSP_170_p;
  assign addKernel_41_A_2 = dSP_298_p;
  assign addKernel_41_A_3 = dSP_426_p;
  assign addKernel_41_A_4 = dSP_554_p;
  assign addKernel_41_A_5 = dSP_682_p;
  assign addKernel_41_A_6 = dSP_810_p;
  assign addKernel_41_A_7 = dSP_938_p;
  assign addKernel_41_A_8 = dSP_1066_p;
  assign addKernel_42_A_0 = dSP_43_p;
  assign addKernel_42_A_1 = dSP_171_p;
  assign addKernel_42_A_2 = dSP_299_p;
  assign addKernel_42_A_3 = dSP_427_p;
  assign addKernel_42_A_4 = dSP_555_p;
  assign addKernel_42_A_5 = dSP_683_p;
  assign addKernel_42_A_6 = dSP_811_p;
  assign addKernel_42_A_7 = dSP_939_p;
  assign addKernel_42_A_8 = dSP_1067_p;
  assign addKernel_43_A_0 = dSP_44_p;
  assign addKernel_43_A_1 = dSP_172_p;
  assign addKernel_43_A_2 = dSP_300_p;
  assign addKernel_43_A_3 = dSP_428_p;
  assign addKernel_43_A_4 = dSP_556_p;
  assign addKernel_43_A_5 = dSP_684_p;
  assign addKernel_43_A_6 = dSP_812_p;
  assign addKernel_43_A_7 = dSP_940_p;
  assign addKernel_43_A_8 = dSP_1068_p;
  assign addKernel_44_A_0 = dSP_45_p;
  assign addKernel_44_A_1 = dSP_173_p;
  assign addKernel_44_A_2 = dSP_301_p;
  assign addKernel_44_A_3 = dSP_429_p;
  assign addKernel_44_A_4 = dSP_557_p;
  assign addKernel_44_A_5 = dSP_685_p;
  assign addKernel_44_A_6 = dSP_813_p;
  assign addKernel_44_A_7 = dSP_941_p;
  assign addKernel_44_A_8 = dSP_1069_p;
  assign addKernel_45_A_0 = dSP_46_p;
  assign addKernel_45_A_1 = dSP_174_p;
  assign addKernel_45_A_2 = dSP_302_p;
  assign addKernel_45_A_3 = dSP_430_p;
  assign addKernel_45_A_4 = dSP_558_p;
  assign addKernel_45_A_5 = dSP_686_p;
  assign addKernel_45_A_6 = dSP_814_p;
  assign addKernel_45_A_7 = dSP_942_p;
  assign addKernel_45_A_8 = dSP_1070_p;
  assign addKernel_46_A_0 = dSP_47_p;
  assign addKernel_46_A_1 = dSP_175_p;
  assign addKernel_46_A_2 = dSP_303_p;
  assign addKernel_46_A_3 = dSP_431_p;
  assign addKernel_46_A_4 = dSP_559_p;
  assign addKernel_46_A_5 = dSP_687_p;
  assign addKernel_46_A_6 = dSP_815_p;
  assign addKernel_46_A_7 = dSP_943_p;
  assign addKernel_46_A_8 = dSP_1071_p;
  assign addKernel_47_A_0 = dSP_48_p;
  assign addKernel_47_A_1 = dSP_176_p;
  assign addKernel_47_A_2 = dSP_304_p;
  assign addKernel_47_A_3 = dSP_432_p;
  assign addKernel_47_A_4 = dSP_560_p;
  assign addKernel_47_A_5 = dSP_688_p;
  assign addKernel_47_A_6 = dSP_816_p;
  assign addKernel_47_A_7 = dSP_944_p;
  assign addKernel_47_A_8 = dSP_1072_p;
  assign addKernel_48_A_0 = dSP_49_p;
  assign addKernel_48_A_1 = dSP_177_p;
  assign addKernel_48_A_2 = dSP_305_p;
  assign addKernel_48_A_3 = dSP_433_p;
  assign addKernel_48_A_4 = dSP_561_p;
  assign addKernel_48_A_5 = dSP_689_p;
  assign addKernel_48_A_6 = dSP_817_p;
  assign addKernel_48_A_7 = dSP_945_p;
  assign addKernel_48_A_8 = dSP_1073_p;
  assign addKernel_49_A_0 = dSP_50_p;
  assign addKernel_49_A_1 = dSP_178_p;
  assign addKernel_49_A_2 = dSP_306_p;
  assign addKernel_49_A_3 = dSP_434_p;
  assign addKernel_49_A_4 = dSP_562_p;
  assign addKernel_49_A_5 = dSP_690_p;
  assign addKernel_49_A_6 = dSP_818_p;
  assign addKernel_49_A_7 = dSP_946_p;
  assign addKernel_49_A_8 = dSP_1074_p;
  assign addKernel_50_A_0 = dSP_51_p;
  assign addKernel_50_A_1 = dSP_179_p;
  assign addKernel_50_A_2 = dSP_307_p;
  assign addKernel_50_A_3 = dSP_435_p;
  assign addKernel_50_A_4 = dSP_563_p;
  assign addKernel_50_A_5 = dSP_691_p;
  assign addKernel_50_A_6 = dSP_819_p;
  assign addKernel_50_A_7 = dSP_947_p;
  assign addKernel_50_A_8 = dSP_1075_p;
  assign addKernel_51_A_0 = dSP_52_p;
  assign addKernel_51_A_1 = dSP_180_p;
  assign addKernel_51_A_2 = dSP_308_p;
  assign addKernel_51_A_3 = dSP_436_p;
  assign addKernel_51_A_4 = dSP_564_p;
  assign addKernel_51_A_5 = dSP_692_p;
  assign addKernel_51_A_6 = dSP_820_p;
  assign addKernel_51_A_7 = dSP_948_p;
  assign addKernel_51_A_8 = dSP_1076_p;
  assign addKernel_52_A_0 = dSP_53_p;
  assign addKernel_52_A_1 = dSP_181_p;
  assign addKernel_52_A_2 = dSP_309_p;
  assign addKernel_52_A_3 = dSP_437_p;
  assign addKernel_52_A_4 = dSP_565_p;
  assign addKernel_52_A_5 = dSP_693_p;
  assign addKernel_52_A_6 = dSP_821_p;
  assign addKernel_52_A_7 = dSP_949_p;
  assign addKernel_52_A_8 = dSP_1077_p;
  assign addKernel_53_A_0 = dSP_54_p;
  assign addKernel_53_A_1 = dSP_182_p;
  assign addKernel_53_A_2 = dSP_310_p;
  assign addKernel_53_A_3 = dSP_438_p;
  assign addKernel_53_A_4 = dSP_566_p;
  assign addKernel_53_A_5 = dSP_694_p;
  assign addKernel_53_A_6 = dSP_822_p;
  assign addKernel_53_A_7 = dSP_950_p;
  assign addKernel_53_A_8 = dSP_1078_p;
  assign addKernel_54_A_0 = dSP_55_p;
  assign addKernel_54_A_1 = dSP_183_p;
  assign addKernel_54_A_2 = dSP_311_p;
  assign addKernel_54_A_3 = dSP_439_p;
  assign addKernel_54_A_4 = dSP_567_p;
  assign addKernel_54_A_5 = dSP_695_p;
  assign addKernel_54_A_6 = dSP_823_p;
  assign addKernel_54_A_7 = dSP_951_p;
  assign addKernel_54_A_8 = dSP_1079_p;
  assign addKernel_55_A_0 = dSP_56_p;
  assign addKernel_55_A_1 = dSP_184_p;
  assign addKernel_55_A_2 = dSP_312_p;
  assign addKernel_55_A_3 = dSP_440_p;
  assign addKernel_55_A_4 = dSP_568_p;
  assign addKernel_55_A_5 = dSP_696_p;
  assign addKernel_55_A_6 = dSP_824_p;
  assign addKernel_55_A_7 = dSP_952_p;
  assign addKernel_55_A_8 = dSP_1080_p;
  assign addKernel_56_A_0 = dSP_57_p;
  assign addKernel_56_A_1 = dSP_185_p;
  assign addKernel_56_A_2 = dSP_313_p;
  assign addKernel_56_A_3 = dSP_441_p;
  assign addKernel_56_A_4 = dSP_569_p;
  assign addKernel_56_A_5 = dSP_697_p;
  assign addKernel_56_A_6 = dSP_825_p;
  assign addKernel_56_A_7 = dSP_953_p;
  assign addKernel_56_A_8 = dSP_1081_p;
  assign addKernel_57_A_0 = dSP_58_p;
  assign addKernel_57_A_1 = dSP_186_p;
  assign addKernel_57_A_2 = dSP_314_p;
  assign addKernel_57_A_3 = dSP_442_p;
  assign addKernel_57_A_4 = dSP_570_p;
  assign addKernel_57_A_5 = dSP_698_p;
  assign addKernel_57_A_6 = dSP_826_p;
  assign addKernel_57_A_7 = dSP_954_p;
  assign addKernel_57_A_8 = dSP_1082_p;
  assign addKernel_58_A_0 = dSP_59_p;
  assign addKernel_58_A_1 = dSP_187_p;
  assign addKernel_58_A_2 = dSP_315_p;
  assign addKernel_58_A_3 = dSP_443_p;
  assign addKernel_58_A_4 = dSP_571_p;
  assign addKernel_58_A_5 = dSP_699_p;
  assign addKernel_58_A_6 = dSP_827_p;
  assign addKernel_58_A_7 = dSP_955_p;
  assign addKernel_58_A_8 = dSP_1083_p;
  assign addKernel_59_A_0 = dSP_60_p;
  assign addKernel_59_A_1 = dSP_188_p;
  assign addKernel_59_A_2 = dSP_316_p;
  assign addKernel_59_A_3 = dSP_444_p;
  assign addKernel_59_A_4 = dSP_572_p;
  assign addKernel_59_A_5 = dSP_700_p;
  assign addKernel_59_A_6 = dSP_828_p;
  assign addKernel_59_A_7 = dSP_956_p;
  assign addKernel_59_A_8 = dSP_1084_p;
  assign addKernel_60_A_0 = dSP_61_p;
  assign addKernel_60_A_1 = dSP_189_p;
  assign addKernel_60_A_2 = dSP_317_p;
  assign addKernel_60_A_3 = dSP_445_p;
  assign addKernel_60_A_4 = dSP_573_p;
  assign addKernel_60_A_5 = dSP_701_p;
  assign addKernel_60_A_6 = dSP_829_p;
  assign addKernel_60_A_7 = dSP_957_p;
  assign addKernel_60_A_8 = dSP_1085_p;
  assign addKernel_61_A_0 = dSP_62_p;
  assign addKernel_61_A_1 = dSP_190_p;
  assign addKernel_61_A_2 = dSP_318_p;
  assign addKernel_61_A_3 = dSP_446_p;
  assign addKernel_61_A_4 = dSP_574_p;
  assign addKernel_61_A_5 = dSP_702_p;
  assign addKernel_61_A_6 = dSP_830_p;
  assign addKernel_61_A_7 = dSP_958_p;
  assign addKernel_61_A_8 = dSP_1086_p;
  assign addKernel_62_A_0 = dSP_63_p;
  assign addKernel_62_A_1 = dSP_191_p;
  assign addKernel_62_A_2 = dSP_319_p;
  assign addKernel_62_A_3 = dSP_447_p;
  assign addKernel_62_A_4 = dSP_575_p;
  assign addKernel_62_A_5 = dSP_703_p;
  assign addKernel_62_A_6 = dSP_831_p;
  assign addKernel_62_A_7 = dSP_959_p;
  assign addKernel_62_A_8 = dSP_1087_p;
  assign addKernel_63_A_0 = dSP_64_p;
  assign addKernel_63_A_1 = dSP_192_p;
  assign addKernel_63_A_2 = dSP_320_p;
  assign addKernel_63_A_3 = dSP_448_p;
  assign addKernel_63_A_4 = dSP_576_p;
  assign addKernel_63_A_5 = dSP_704_p;
  assign addKernel_63_A_6 = dSP_832_p;
  assign addKernel_63_A_7 = dSP_960_p;
  assign addKernel_63_A_8 = dSP_1088_p;
  assign addKernel_64_A_0 = dSP_65_p;
  assign addKernel_64_A_1 = dSP_193_p;
  assign addKernel_64_A_2 = dSP_321_p;
  assign addKernel_64_A_3 = dSP_449_p;
  assign addKernel_64_A_4 = dSP_577_p;
  assign addKernel_64_A_5 = dSP_705_p;
  assign addKernel_64_A_6 = dSP_833_p;
  assign addKernel_64_A_7 = dSP_961_p;
  assign addKernel_64_A_8 = dSP_1089_p;
  assign addKernel_65_A_0 = dSP_66_p;
  assign addKernel_65_A_1 = dSP_194_p;
  assign addKernel_65_A_2 = dSP_322_p;
  assign addKernel_65_A_3 = dSP_450_p;
  assign addKernel_65_A_4 = dSP_578_p;
  assign addKernel_65_A_5 = dSP_706_p;
  assign addKernel_65_A_6 = dSP_834_p;
  assign addKernel_65_A_7 = dSP_962_p;
  assign addKernel_65_A_8 = dSP_1090_p;
  assign addKernel_66_A_0 = dSP_67_p;
  assign addKernel_66_A_1 = dSP_195_p;
  assign addKernel_66_A_2 = dSP_323_p;
  assign addKernel_66_A_3 = dSP_451_p;
  assign addKernel_66_A_4 = dSP_579_p;
  assign addKernel_66_A_5 = dSP_707_p;
  assign addKernel_66_A_6 = dSP_835_p;
  assign addKernel_66_A_7 = dSP_963_p;
  assign addKernel_66_A_8 = dSP_1091_p;
  assign addKernel_67_A_0 = dSP_68_p;
  assign addKernel_67_A_1 = dSP_196_p;
  assign addKernel_67_A_2 = dSP_324_p;
  assign addKernel_67_A_3 = dSP_452_p;
  assign addKernel_67_A_4 = dSP_580_p;
  assign addKernel_67_A_5 = dSP_708_p;
  assign addKernel_67_A_6 = dSP_836_p;
  assign addKernel_67_A_7 = dSP_964_p;
  assign addKernel_67_A_8 = dSP_1092_p;
  assign addKernel_68_A_0 = dSP_69_p;
  assign addKernel_68_A_1 = dSP_197_p;
  assign addKernel_68_A_2 = dSP_325_p;
  assign addKernel_68_A_3 = dSP_453_p;
  assign addKernel_68_A_4 = dSP_581_p;
  assign addKernel_68_A_5 = dSP_709_p;
  assign addKernel_68_A_6 = dSP_837_p;
  assign addKernel_68_A_7 = dSP_965_p;
  assign addKernel_68_A_8 = dSP_1093_p;
  assign addKernel_69_A_0 = dSP_70_p;
  assign addKernel_69_A_1 = dSP_198_p;
  assign addKernel_69_A_2 = dSP_326_p;
  assign addKernel_69_A_3 = dSP_454_p;
  assign addKernel_69_A_4 = dSP_582_p;
  assign addKernel_69_A_5 = dSP_710_p;
  assign addKernel_69_A_6 = dSP_838_p;
  assign addKernel_69_A_7 = dSP_966_p;
  assign addKernel_69_A_8 = dSP_1094_p;
  assign addKernel_70_A_0 = dSP_71_p;
  assign addKernel_70_A_1 = dSP_199_p;
  assign addKernel_70_A_2 = dSP_327_p;
  assign addKernel_70_A_3 = dSP_455_p;
  assign addKernel_70_A_4 = dSP_583_p;
  assign addKernel_70_A_5 = dSP_711_p;
  assign addKernel_70_A_6 = dSP_839_p;
  assign addKernel_70_A_7 = dSP_967_p;
  assign addKernel_70_A_8 = dSP_1095_p;
  assign addKernel_71_A_0 = dSP_72_p;
  assign addKernel_71_A_1 = dSP_200_p;
  assign addKernel_71_A_2 = dSP_328_p;
  assign addKernel_71_A_3 = dSP_456_p;
  assign addKernel_71_A_4 = dSP_584_p;
  assign addKernel_71_A_5 = dSP_712_p;
  assign addKernel_71_A_6 = dSP_840_p;
  assign addKernel_71_A_7 = dSP_968_p;
  assign addKernel_71_A_8 = dSP_1096_p;
  assign addKernel_72_A_0 = dSP_73_p;
  assign addKernel_72_A_1 = dSP_201_p;
  assign addKernel_72_A_2 = dSP_329_p;
  assign addKernel_72_A_3 = dSP_457_p;
  assign addKernel_72_A_4 = dSP_585_p;
  assign addKernel_72_A_5 = dSP_713_p;
  assign addKernel_72_A_6 = dSP_841_p;
  assign addKernel_72_A_7 = dSP_969_p;
  assign addKernel_72_A_8 = dSP_1097_p;
  assign addKernel_73_A_0 = dSP_74_p;
  assign addKernel_73_A_1 = dSP_202_p;
  assign addKernel_73_A_2 = dSP_330_p;
  assign addKernel_73_A_3 = dSP_458_p;
  assign addKernel_73_A_4 = dSP_586_p;
  assign addKernel_73_A_5 = dSP_714_p;
  assign addKernel_73_A_6 = dSP_842_p;
  assign addKernel_73_A_7 = dSP_970_p;
  assign addKernel_73_A_8 = dSP_1098_p;
  assign addKernel_74_A_0 = dSP_75_p;
  assign addKernel_74_A_1 = dSP_203_p;
  assign addKernel_74_A_2 = dSP_331_p;
  assign addKernel_74_A_3 = dSP_459_p;
  assign addKernel_74_A_4 = dSP_587_p;
  assign addKernel_74_A_5 = dSP_715_p;
  assign addKernel_74_A_6 = dSP_843_p;
  assign addKernel_74_A_7 = dSP_971_p;
  assign addKernel_74_A_8 = dSP_1099_p;
  assign addKernel_75_A_0 = dSP_76_p;
  assign addKernel_75_A_1 = dSP_204_p;
  assign addKernel_75_A_2 = dSP_332_p;
  assign addKernel_75_A_3 = dSP_460_p;
  assign addKernel_75_A_4 = dSP_588_p;
  assign addKernel_75_A_5 = dSP_716_p;
  assign addKernel_75_A_6 = dSP_844_p;
  assign addKernel_75_A_7 = dSP_972_p;
  assign addKernel_75_A_8 = dSP_1100_p;
  assign addKernel_76_A_0 = dSP_77_p;
  assign addKernel_76_A_1 = dSP_205_p;
  assign addKernel_76_A_2 = dSP_333_p;
  assign addKernel_76_A_3 = dSP_461_p;
  assign addKernel_76_A_4 = dSP_589_p;
  assign addKernel_76_A_5 = dSP_717_p;
  assign addKernel_76_A_6 = dSP_845_p;
  assign addKernel_76_A_7 = dSP_973_p;
  assign addKernel_76_A_8 = dSP_1101_p;
  assign addKernel_77_A_0 = dSP_78_p;
  assign addKernel_77_A_1 = dSP_206_p;
  assign addKernel_77_A_2 = dSP_334_p;
  assign addKernel_77_A_3 = dSP_462_p;
  assign addKernel_77_A_4 = dSP_590_p;
  assign addKernel_77_A_5 = dSP_718_p;
  assign addKernel_77_A_6 = dSP_846_p;
  assign addKernel_77_A_7 = dSP_974_p;
  assign addKernel_77_A_8 = dSP_1102_p;
  assign addKernel_78_A_0 = dSP_79_p;
  assign addKernel_78_A_1 = dSP_207_p;
  assign addKernel_78_A_2 = dSP_335_p;
  assign addKernel_78_A_3 = dSP_463_p;
  assign addKernel_78_A_4 = dSP_591_p;
  assign addKernel_78_A_5 = dSP_719_p;
  assign addKernel_78_A_6 = dSP_847_p;
  assign addKernel_78_A_7 = dSP_975_p;
  assign addKernel_78_A_8 = dSP_1103_p;
  assign addKernel_79_A_0 = dSP_80_p;
  assign addKernel_79_A_1 = dSP_208_p;
  assign addKernel_79_A_2 = dSP_336_p;
  assign addKernel_79_A_3 = dSP_464_p;
  assign addKernel_79_A_4 = dSP_592_p;
  assign addKernel_79_A_5 = dSP_720_p;
  assign addKernel_79_A_6 = dSP_848_p;
  assign addKernel_79_A_7 = dSP_976_p;
  assign addKernel_79_A_8 = dSP_1104_p;
  assign addKernel_80_A_0 = dSP_81_p;
  assign addKernel_80_A_1 = dSP_209_p;
  assign addKernel_80_A_2 = dSP_337_p;
  assign addKernel_80_A_3 = dSP_465_p;
  assign addKernel_80_A_4 = dSP_593_p;
  assign addKernel_80_A_5 = dSP_721_p;
  assign addKernel_80_A_6 = dSP_849_p;
  assign addKernel_80_A_7 = dSP_977_p;
  assign addKernel_80_A_8 = dSP_1105_p;
  assign addKernel_81_A_0 = dSP_82_p;
  assign addKernel_81_A_1 = dSP_210_p;
  assign addKernel_81_A_2 = dSP_338_p;
  assign addKernel_81_A_3 = dSP_466_p;
  assign addKernel_81_A_4 = dSP_594_p;
  assign addKernel_81_A_5 = dSP_722_p;
  assign addKernel_81_A_6 = dSP_850_p;
  assign addKernel_81_A_7 = dSP_978_p;
  assign addKernel_81_A_8 = dSP_1106_p;
  assign addKernel_82_A_0 = dSP_83_p;
  assign addKernel_82_A_1 = dSP_211_p;
  assign addKernel_82_A_2 = dSP_339_p;
  assign addKernel_82_A_3 = dSP_467_p;
  assign addKernel_82_A_4 = dSP_595_p;
  assign addKernel_82_A_5 = dSP_723_p;
  assign addKernel_82_A_6 = dSP_851_p;
  assign addKernel_82_A_7 = dSP_979_p;
  assign addKernel_82_A_8 = dSP_1107_p;
  assign addKernel_83_A_0 = dSP_84_p;
  assign addKernel_83_A_1 = dSP_212_p;
  assign addKernel_83_A_2 = dSP_340_p;
  assign addKernel_83_A_3 = dSP_468_p;
  assign addKernel_83_A_4 = dSP_596_p;
  assign addKernel_83_A_5 = dSP_724_p;
  assign addKernel_83_A_6 = dSP_852_p;
  assign addKernel_83_A_7 = dSP_980_p;
  assign addKernel_83_A_8 = dSP_1108_p;
  assign addKernel_84_A_0 = dSP_85_p;
  assign addKernel_84_A_1 = dSP_213_p;
  assign addKernel_84_A_2 = dSP_341_p;
  assign addKernel_84_A_3 = dSP_469_p;
  assign addKernel_84_A_4 = dSP_597_p;
  assign addKernel_84_A_5 = dSP_725_p;
  assign addKernel_84_A_6 = dSP_853_p;
  assign addKernel_84_A_7 = dSP_981_p;
  assign addKernel_84_A_8 = dSP_1109_p;
  assign addKernel_85_A_0 = dSP_86_p;
  assign addKernel_85_A_1 = dSP_214_p;
  assign addKernel_85_A_2 = dSP_342_p;
  assign addKernel_85_A_3 = dSP_470_p;
  assign addKernel_85_A_4 = dSP_598_p;
  assign addKernel_85_A_5 = dSP_726_p;
  assign addKernel_85_A_6 = dSP_854_p;
  assign addKernel_85_A_7 = dSP_982_p;
  assign addKernel_85_A_8 = dSP_1110_p;
  assign addKernel_86_A_0 = dSP_87_p;
  assign addKernel_86_A_1 = dSP_215_p;
  assign addKernel_86_A_2 = dSP_343_p;
  assign addKernel_86_A_3 = dSP_471_p;
  assign addKernel_86_A_4 = dSP_599_p;
  assign addKernel_86_A_5 = dSP_727_p;
  assign addKernel_86_A_6 = dSP_855_p;
  assign addKernel_86_A_7 = dSP_983_p;
  assign addKernel_86_A_8 = dSP_1111_p;
  assign addKernel_87_A_0 = dSP_88_p;
  assign addKernel_87_A_1 = dSP_216_p;
  assign addKernel_87_A_2 = dSP_344_p;
  assign addKernel_87_A_3 = dSP_472_p;
  assign addKernel_87_A_4 = dSP_600_p;
  assign addKernel_87_A_5 = dSP_728_p;
  assign addKernel_87_A_6 = dSP_856_p;
  assign addKernel_87_A_7 = dSP_984_p;
  assign addKernel_87_A_8 = dSP_1112_p;
  assign addKernel_88_A_0 = dSP_89_p;
  assign addKernel_88_A_1 = dSP_217_p;
  assign addKernel_88_A_2 = dSP_345_p;
  assign addKernel_88_A_3 = dSP_473_p;
  assign addKernel_88_A_4 = dSP_601_p;
  assign addKernel_88_A_5 = dSP_729_p;
  assign addKernel_88_A_6 = dSP_857_p;
  assign addKernel_88_A_7 = dSP_985_p;
  assign addKernel_88_A_8 = dSP_1113_p;
  assign addKernel_89_A_0 = dSP_90_p;
  assign addKernel_89_A_1 = dSP_218_p;
  assign addKernel_89_A_2 = dSP_346_p;
  assign addKernel_89_A_3 = dSP_474_p;
  assign addKernel_89_A_4 = dSP_602_p;
  assign addKernel_89_A_5 = dSP_730_p;
  assign addKernel_89_A_6 = dSP_858_p;
  assign addKernel_89_A_7 = dSP_986_p;
  assign addKernel_89_A_8 = dSP_1114_p;
  assign addKernel_90_A_0 = dSP_91_p;
  assign addKernel_90_A_1 = dSP_219_p;
  assign addKernel_90_A_2 = dSP_347_p;
  assign addKernel_90_A_3 = dSP_475_p;
  assign addKernel_90_A_4 = dSP_603_p;
  assign addKernel_90_A_5 = dSP_731_p;
  assign addKernel_90_A_6 = dSP_859_p;
  assign addKernel_90_A_7 = dSP_987_p;
  assign addKernel_90_A_8 = dSP_1115_p;
  assign addKernel_91_A_0 = dSP_92_p;
  assign addKernel_91_A_1 = dSP_220_p;
  assign addKernel_91_A_2 = dSP_348_p;
  assign addKernel_91_A_3 = dSP_476_p;
  assign addKernel_91_A_4 = dSP_604_p;
  assign addKernel_91_A_5 = dSP_732_p;
  assign addKernel_91_A_6 = dSP_860_p;
  assign addKernel_91_A_7 = dSP_988_p;
  assign addKernel_91_A_8 = dSP_1116_p;
  assign addKernel_92_A_0 = dSP_93_p;
  assign addKernel_92_A_1 = dSP_221_p;
  assign addKernel_92_A_2 = dSP_349_p;
  assign addKernel_92_A_3 = dSP_477_p;
  assign addKernel_92_A_4 = dSP_605_p;
  assign addKernel_92_A_5 = dSP_733_p;
  assign addKernel_92_A_6 = dSP_861_p;
  assign addKernel_92_A_7 = dSP_989_p;
  assign addKernel_92_A_8 = dSP_1117_p;
  assign addKernel_93_A_0 = dSP_94_p;
  assign addKernel_93_A_1 = dSP_222_p;
  assign addKernel_93_A_2 = dSP_350_p;
  assign addKernel_93_A_3 = dSP_478_p;
  assign addKernel_93_A_4 = dSP_606_p;
  assign addKernel_93_A_5 = dSP_734_p;
  assign addKernel_93_A_6 = dSP_862_p;
  assign addKernel_93_A_7 = dSP_990_p;
  assign addKernel_93_A_8 = dSP_1118_p;
  assign addKernel_94_A_0 = dSP_95_p;
  assign addKernel_94_A_1 = dSP_223_p;
  assign addKernel_94_A_2 = dSP_351_p;
  assign addKernel_94_A_3 = dSP_479_p;
  assign addKernel_94_A_4 = dSP_607_p;
  assign addKernel_94_A_5 = dSP_735_p;
  assign addKernel_94_A_6 = dSP_863_p;
  assign addKernel_94_A_7 = dSP_991_p;
  assign addKernel_94_A_8 = dSP_1119_p;
  assign addKernel_95_A_0 = dSP_96_p;
  assign addKernel_95_A_1 = dSP_224_p;
  assign addKernel_95_A_2 = dSP_352_p;
  assign addKernel_95_A_3 = dSP_480_p;
  assign addKernel_95_A_4 = dSP_608_p;
  assign addKernel_95_A_5 = dSP_736_p;
  assign addKernel_95_A_6 = dSP_864_p;
  assign addKernel_95_A_7 = dSP_992_p;
  assign addKernel_95_A_8 = dSP_1120_p;
  assign addKernel_96_A_0 = dSP_97_p;
  assign addKernel_96_A_1 = dSP_225_p;
  assign addKernel_96_A_2 = dSP_353_p;
  assign addKernel_96_A_3 = dSP_481_p;
  assign addKernel_96_A_4 = dSP_609_p;
  assign addKernel_96_A_5 = dSP_737_p;
  assign addKernel_96_A_6 = dSP_865_p;
  assign addKernel_96_A_7 = dSP_993_p;
  assign addKernel_96_A_8 = dSP_1121_p;
  assign addKernel_97_A_0 = dSP_98_p;
  assign addKernel_97_A_1 = dSP_226_p;
  assign addKernel_97_A_2 = dSP_354_p;
  assign addKernel_97_A_3 = dSP_482_p;
  assign addKernel_97_A_4 = dSP_610_p;
  assign addKernel_97_A_5 = dSP_738_p;
  assign addKernel_97_A_6 = dSP_866_p;
  assign addKernel_97_A_7 = dSP_994_p;
  assign addKernel_97_A_8 = dSP_1122_p;
  assign addKernel_98_A_0 = dSP_99_p;
  assign addKernel_98_A_1 = dSP_227_p;
  assign addKernel_98_A_2 = dSP_355_p;
  assign addKernel_98_A_3 = dSP_483_p;
  assign addKernel_98_A_4 = dSP_611_p;
  assign addKernel_98_A_5 = dSP_739_p;
  assign addKernel_98_A_6 = dSP_867_p;
  assign addKernel_98_A_7 = dSP_995_p;
  assign addKernel_98_A_8 = dSP_1123_p;
  assign addKernel_99_A_0 = dSP_100_p;
  assign addKernel_99_A_1 = dSP_228_p;
  assign addKernel_99_A_2 = dSP_356_p;
  assign addKernel_99_A_3 = dSP_484_p;
  assign addKernel_99_A_4 = dSP_612_p;
  assign addKernel_99_A_5 = dSP_740_p;
  assign addKernel_99_A_6 = dSP_868_p;
  assign addKernel_99_A_7 = dSP_996_p;
  assign addKernel_99_A_8 = dSP_1124_p;
  assign addKernel_100_A_0 = dSP_101_p;
  assign addKernel_100_A_1 = dSP_229_p;
  assign addKernel_100_A_2 = dSP_357_p;
  assign addKernel_100_A_3 = dSP_485_p;
  assign addKernel_100_A_4 = dSP_613_p;
  assign addKernel_100_A_5 = dSP_741_p;
  assign addKernel_100_A_6 = dSP_869_p;
  assign addKernel_100_A_7 = dSP_997_p;
  assign addKernel_100_A_8 = dSP_1125_p;
  assign addKernel_101_A_0 = dSP_102_p;
  assign addKernel_101_A_1 = dSP_230_p;
  assign addKernel_101_A_2 = dSP_358_p;
  assign addKernel_101_A_3 = dSP_486_p;
  assign addKernel_101_A_4 = dSP_614_p;
  assign addKernel_101_A_5 = dSP_742_p;
  assign addKernel_101_A_6 = dSP_870_p;
  assign addKernel_101_A_7 = dSP_998_p;
  assign addKernel_101_A_8 = dSP_1126_p;
  assign addKernel_102_A_0 = dSP_103_p;
  assign addKernel_102_A_1 = dSP_231_p;
  assign addKernel_102_A_2 = dSP_359_p;
  assign addKernel_102_A_3 = dSP_487_p;
  assign addKernel_102_A_4 = dSP_615_p;
  assign addKernel_102_A_5 = dSP_743_p;
  assign addKernel_102_A_6 = dSP_871_p;
  assign addKernel_102_A_7 = dSP_999_p;
  assign addKernel_102_A_8 = dSP_1127_p;
  assign addKernel_103_A_0 = dSP_104_p;
  assign addKernel_103_A_1 = dSP_232_p;
  assign addKernel_103_A_2 = dSP_360_p;
  assign addKernel_103_A_3 = dSP_488_p;
  assign addKernel_103_A_4 = dSP_616_p;
  assign addKernel_103_A_5 = dSP_744_p;
  assign addKernel_103_A_6 = dSP_872_p;
  assign addKernel_103_A_7 = dSP_1000_p;
  assign addKernel_103_A_8 = dSP_1128_p;
  assign addKernel_104_A_0 = dSP_105_p;
  assign addKernel_104_A_1 = dSP_233_p;
  assign addKernel_104_A_2 = dSP_361_p;
  assign addKernel_104_A_3 = dSP_489_p;
  assign addKernel_104_A_4 = dSP_617_p;
  assign addKernel_104_A_5 = dSP_745_p;
  assign addKernel_104_A_6 = dSP_873_p;
  assign addKernel_104_A_7 = dSP_1001_p;
  assign addKernel_104_A_8 = dSP_1129_p;
  assign addKernel_105_A_0 = dSP_106_p;
  assign addKernel_105_A_1 = dSP_234_p;
  assign addKernel_105_A_2 = dSP_362_p;
  assign addKernel_105_A_3 = dSP_490_p;
  assign addKernel_105_A_4 = dSP_618_p;
  assign addKernel_105_A_5 = dSP_746_p;
  assign addKernel_105_A_6 = dSP_874_p;
  assign addKernel_105_A_7 = dSP_1002_p;
  assign addKernel_105_A_8 = dSP_1130_p;
  assign addKernel_106_A_0 = dSP_107_p;
  assign addKernel_106_A_1 = dSP_235_p;
  assign addKernel_106_A_2 = dSP_363_p;
  assign addKernel_106_A_3 = dSP_491_p;
  assign addKernel_106_A_4 = dSP_619_p;
  assign addKernel_106_A_5 = dSP_747_p;
  assign addKernel_106_A_6 = dSP_875_p;
  assign addKernel_106_A_7 = dSP_1003_p;
  assign addKernel_106_A_8 = dSP_1131_p;
  assign addKernel_107_A_0 = dSP_108_p;
  assign addKernel_107_A_1 = dSP_236_p;
  assign addKernel_107_A_2 = dSP_364_p;
  assign addKernel_107_A_3 = dSP_492_p;
  assign addKernel_107_A_4 = dSP_620_p;
  assign addKernel_107_A_5 = dSP_748_p;
  assign addKernel_107_A_6 = dSP_876_p;
  assign addKernel_107_A_7 = dSP_1004_p;
  assign addKernel_107_A_8 = dSP_1132_p;
  assign addKernel_108_A_0 = dSP_109_p;
  assign addKernel_108_A_1 = dSP_237_p;
  assign addKernel_108_A_2 = dSP_365_p;
  assign addKernel_108_A_3 = dSP_493_p;
  assign addKernel_108_A_4 = dSP_621_p;
  assign addKernel_108_A_5 = dSP_749_p;
  assign addKernel_108_A_6 = dSP_877_p;
  assign addKernel_108_A_7 = dSP_1005_p;
  assign addKernel_108_A_8 = dSP_1133_p;
  assign addKernel_109_A_0 = dSP_110_p;
  assign addKernel_109_A_1 = dSP_238_p;
  assign addKernel_109_A_2 = dSP_366_p;
  assign addKernel_109_A_3 = dSP_494_p;
  assign addKernel_109_A_4 = dSP_622_p;
  assign addKernel_109_A_5 = dSP_750_p;
  assign addKernel_109_A_6 = dSP_878_p;
  assign addKernel_109_A_7 = dSP_1006_p;
  assign addKernel_109_A_8 = dSP_1134_p;
  assign addKernel_110_A_0 = dSP_111_p;
  assign addKernel_110_A_1 = dSP_239_p;
  assign addKernel_110_A_2 = dSP_367_p;
  assign addKernel_110_A_3 = dSP_495_p;
  assign addKernel_110_A_4 = dSP_623_p;
  assign addKernel_110_A_5 = dSP_751_p;
  assign addKernel_110_A_6 = dSP_879_p;
  assign addKernel_110_A_7 = dSP_1007_p;
  assign addKernel_110_A_8 = dSP_1135_p;
  assign addKernel_111_A_0 = dSP_112_p;
  assign addKernel_111_A_1 = dSP_240_p;
  assign addKernel_111_A_2 = dSP_368_p;
  assign addKernel_111_A_3 = dSP_496_p;
  assign addKernel_111_A_4 = dSP_624_p;
  assign addKernel_111_A_5 = dSP_752_p;
  assign addKernel_111_A_6 = dSP_880_p;
  assign addKernel_111_A_7 = dSP_1008_p;
  assign addKernel_111_A_8 = dSP_1136_p;
  assign addKernel_112_A_0 = dSP_113_p;
  assign addKernel_112_A_1 = dSP_241_p;
  assign addKernel_112_A_2 = dSP_369_p;
  assign addKernel_112_A_3 = dSP_497_p;
  assign addKernel_112_A_4 = dSP_625_p;
  assign addKernel_112_A_5 = dSP_753_p;
  assign addKernel_112_A_6 = dSP_881_p;
  assign addKernel_112_A_7 = dSP_1009_p;
  assign addKernel_112_A_8 = dSP_1137_p;
  assign addKernel_113_A_0 = dSP_114_p;
  assign addKernel_113_A_1 = dSP_242_p;
  assign addKernel_113_A_2 = dSP_370_p;
  assign addKernel_113_A_3 = dSP_498_p;
  assign addKernel_113_A_4 = dSP_626_p;
  assign addKernel_113_A_5 = dSP_754_p;
  assign addKernel_113_A_6 = dSP_882_p;
  assign addKernel_113_A_7 = dSP_1010_p;
  assign addKernel_113_A_8 = dSP_1138_p;
  assign addKernel_114_A_0 = dSP_115_p;
  assign addKernel_114_A_1 = dSP_243_p;
  assign addKernel_114_A_2 = dSP_371_p;
  assign addKernel_114_A_3 = dSP_499_p;
  assign addKernel_114_A_4 = dSP_627_p;
  assign addKernel_114_A_5 = dSP_755_p;
  assign addKernel_114_A_6 = dSP_883_p;
  assign addKernel_114_A_7 = dSP_1011_p;
  assign addKernel_114_A_8 = dSP_1139_p;
  assign addKernel_115_A_0 = dSP_116_p;
  assign addKernel_115_A_1 = dSP_244_p;
  assign addKernel_115_A_2 = dSP_372_p;
  assign addKernel_115_A_3 = dSP_500_p;
  assign addKernel_115_A_4 = dSP_628_p;
  assign addKernel_115_A_5 = dSP_756_p;
  assign addKernel_115_A_6 = dSP_884_p;
  assign addKernel_115_A_7 = dSP_1012_p;
  assign addKernel_115_A_8 = dSP_1140_p;
  assign addKernel_116_A_0 = dSP_117_p;
  assign addKernel_116_A_1 = dSP_245_p;
  assign addKernel_116_A_2 = dSP_373_p;
  assign addKernel_116_A_3 = dSP_501_p;
  assign addKernel_116_A_4 = dSP_629_p;
  assign addKernel_116_A_5 = dSP_757_p;
  assign addKernel_116_A_6 = dSP_885_p;
  assign addKernel_116_A_7 = dSP_1013_p;
  assign addKernel_116_A_8 = dSP_1141_p;
  assign addKernel_117_A_0 = dSP_118_p;
  assign addKernel_117_A_1 = dSP_246_p;
  assign addKernel_117_A_2 = dSP_374_p;
  assign addKernel_117_A_3 = dSP_502_p;
  assign addKernel_117_A_4 = dSP_630_p;
  assign addKernel_117_A_5 = dSP_758_p;
  assign addKernel_117_A_6 = dSP_886_p;
  assign addKernel_117_A_7 = dSP_1014_p;
  assign addKernel_117_A_8 = dSP_1142_p;
  assign addKernel_118_A_0 = dSP_119_p;
  assign addKernel_118_A_1 = dSP_247_p;
  assign addKernel_118_A_2 = dSP_375_p;
  assign addKernel_118_A_3 = dSP_503_p;
  assign addKernel_118_A_4 = dSP_631_p;
  assign addKernel_118_A_5 = dSP_759_p;
  assign addKernel_118_A_6 = dSP_887_p;
  assign addKernel_118_A_7 = dSP_1015_p;
  assign addKernel_118_A_8 = dSP_1143_p;
  assign addKernel_119_A_0 = dSP_120_p;
  assign addKernel_119_A_1 = dSP_248_p;
  assign addKernel_119_A_2 = dSP_376_p;
  assign addKernel_119_A_3 = dSP_504_p;
  assign addKernel_119_A_4 = dSP_632_p;
  assign addKernel_119_A_5 = dSP_760_p;
  assign addKernel_119_A_6 = dSP_888_p;
  assign addKernel_119_A_7 = dSP_1016_p;
  assign addKernel_119_A_8 = dSP_1144_p;
  assign addKernel_120_A_0 = dSP_121_p;
  assign addKernel_120_A_1 = dSP_249_p;
  assign addKernel_120_A_2 = dSP_377_p;
  assign addKernel_120_A_3 = dSP_505_p;
  assign addKernel_120_A_4 = dSP_633_p;
  assign addKernel_120_A_5 = dSP_761_p;
  assign addKernel_120_A_6 = dSP_889_p;
  assign addKernel_120_A_7 = dSP_1017_p;
  assign addKernel_120_A_8 = dSP_1145_p;
  assign addKernel_121_A_0 = dSP_122_p;
  assign addKernel_121_A_1 = dSP_250_p;
  assign addKernel_121_A_2 = dSP_378_p;
  assign addKernel_121_A_3 = dSP_506_p;
  assign addKernel_121_A_4 = dSP_634_p;
  assign addKernel_121_A_5 = dSP_762_p;
  assign addKernel_121_A_6 = dSP_890_p;
  assign addKernel_121_A_7 = dSP_1018_p;
  assign addKernel_121_A_8 = dSP_1146_p;
  assign addKernel_122_A_0 = dSP_123_p;
  assign addKernel_122_A_1 = dSP_251_p;
  assign addKernel_122_A_2 = dSP_379_p;
  assign addKernel_122_A_3 = dSP_507_p;
  assign addKernel_122_A_4 = dSP_635_p;
  assign addKernel_122_A_5 = dSP_763_p;
  assign addKernel_122_A_6 = dSP_891_p;
  assign addKernel_122_A_7 = dSP_1019_p;
  assign addKernel_122_A_8 = dSP_1147_p;
  assign addKernel_123_A_0 = dSP_124_p;
  assign addKernel_123_A_1 = dSP_252_p;
  assign addKernel_123_A_2 = dSP_380_p;
  assign addKernel_123_A_3 = dSP_508_p;
  assign addKernel_123_A_4 = dSP_636_p;
  assign addKernel_123_A_5 = dSP_764_p;
  assign addKernel_123_A_6 = dSP_892_p;
  assign addKernel_123_A_7 = dSP_1020_p;
  assign addKernel_123_A_8 = dSP_1148_p;
  assign addKernel_124_A_0 = dSP_125_p;
  assign addKernel_124_A_1 = dSP_253_p;
  assign addKernel_124_A_2 = dSP_381_p;
  assign addKernel_124_A_3 = dSP_509_p;
  assign addKernel_124_A_4 = dSP_637_p;
  assign addKernel_124_A_5 = dSP_765_p;
  assign addKernel_124_A_6 = dSP_893_p;
  assign addKernel_124_A_7 = dSP_1021_p;
  assign addKernel_124_A_8 = dSP_1149_p;
  assign addKernel_125_A_0 = dSP_126_p;
  assign addKernel_125_A_1 = dSP_254_p;
  assign addKernel_125_A_2 = dSP_382_p;
  assign addKernel_125_A_3 = dSP_510_p;
  assign addKernel_125_A_4 = dSP_638_p;
  assign addKernel_125_A_5 = dSP_766_p;
  assign addKernel_125_A_6 = dSP_894_p;
  assign addKernel_125_A_7 = dSP_1022_p;
  assign addKernel_125_A_8 = dSP_1150_p;
  assign addKernel_126_A_0 = dSP_127_p;
  assign addKernel_126_A_1 = dSP_255_p;
  assign addKernel_126_A_2 = dSP_383_p;
  assign addKernel_126_A_3 = dSP_511_p;
  assign addKernel_126_A_4 = dSP_639_p;
  assign addKernel_126_A_5 = dSP_767_p;
  assign addKernel_126_A_6 = dSP_895_p;
  assign addKernel_126_A_7 = dSP_1023_p;
  assign addKernel_126_A_8 = dSP_1151_p;
  assign addKernel_127_A_0 = dSP_128_p;
  assign addKernel_127_A_1 = dSP_256_p;
  assign addKernel_127_A_2 = dSP_384_p;
  assign addKernel_127_A_3 = dSP_512_p;
  assign addKernel_127_A_4 = dSP_640_p;
  assign addKernel_127_A_5 = dSP_768_p;
  assign addKernel_127_A_6 = dSP_896_p;
  assign addKernel_127_A_7 = dSP_1024_p;
  assign addKernel_127_A_8 = dSP_1152_p;
  assign _zz_A = xAddTimes_136_S;
  assign _zz_A_1 = xAddTimes_137_S;
  assign _zz_A_2 = xAddTimes_138_S;
  assign _zz_A_3 = xAddTimes_139_S;
  assign _zz_A_4 = xAddTimes_140_S;
  assign _zz_A_5 = xAddTimes_141_S;
  assign _zz_A_6 = xAddTimes_142_S;
  assign _zz_A_7 = xAddTimes_143_S;
  assign xAddChannelTimes_16_A = _zz_A[23 : 0];
  assign xAddChannelTimes_17_A = _zz_A[47 : 24];
  assign xAddChannelTimes_18_A = _zz_A_1[23 : 0];
  assign xAddChannelTimes_19_A = _zz_A_1[47 : 24];
  assign xAddChannelTimes_20_A = _zz_A_2[23 : 0];
  assign xAddChannelTimes_21_A = _zz_A_2[47 : 24];
  assign xAddChannelTimes_22_A = _zz_A_3[23 : 0];
  assign xAddChannelTimes_23_A = _zz_A_3[47 : 24];
  assign xAddChannelTimes_24_A = _zz_A_4[23 : 0];
  assign xAddChannelTimes_25_A = _zz_A_4[47 : 24];
  assign xAddChannelTimes_26_A = _zz_A_5[23 : 0];
  assign xAddChannelTimes_27_A = _zz_A_5[47 : 24];
  assign xAddChannelTimes_28_A = _zz_A_6[23 : 0];
  assign xAddChannelTimes_29_A = _zz_A_6[47 : 24];
  assign xAddChannelTimes_30_A = _zz_A_7[23 : 0];
  assign xAddChannelTimes_31_A = _zz_A_7[47 : 24];
  assign mFeatureData_valid = stride_1_mData_valid;
  assign mFeatureData_payload = stride_1_mData_payload;
  assign computeComplete = stride_1_complete;
  assign last = stride_1_last;
  always @(posedge clk) begin
    if(startPa) begin
      _zz_convType <= convType;
    end
    _zz_b_9 <= _zz__zz_1_port1;
    _zz_b_10 <= _zz_b_9;
    _zz_b_11 <= _zz_b_10;
    _zz_b_12 <= _zz_b_11;
    _zz_b_13 <= _zz_b_12;
    _zz_b_14 <= _zz_b_13;
    _zz_b_15 <= _zz_b_14;
    _zz_b_16 <= _zz_b_15;
    _zz_b_17 <= _zz_b_16;
    _zz_b_18 <= _zz_b_17;
    _zz_b_19 <= _zz__zz_2_port1;
    _zz_b_20 <= _zz_b_19;
    _zz_b_21 <= _zz_b_20;
    _zz_b_22 <= _zz_b_21;
    _zz_b_23 <= _zz_b_22;
    _zz_b_24 <= _zz_b_23;
    _zz_b_25 <= _zz_b_24;
    _zz_b_26 <= _zz_b_25;
    _zz_b_27 <= _zz_b_26;
    _zz_b_28 <= _zz_b_27;
    _zz_b_29 <= _zz__zz_3_port1;
    _zz_b_30 <= _zz_b_29;
    _zz_b_31 <= _zz_b_30;
    _zz_b_32 <= _zz_b_31;
    _zz_b_33 <= _zz_b_32;
    _zz_b_34 <= _zz_b_33;
    _zz_b_35 <= _zz_b_34;
    _zz_b_36 <= _zz_b_35;
    _zz_b_37 <= _zz_b_36;
    _zz_b_38 <= _zz_b_37;
    _zz_b_39 <= _zz__zz_4_port1;
    _zz_b_40 <= _zz_b_39;
    _zz_b_41 <= _zz_b_40;
    _zz_b_42 <= _zz_b_41;
    _zz_b_43 <= _zz_b_42;
    _zz_b_44 <= _zz_b_43;
    _zz_b_45 <= _zz_b_44;
    _zz_b_46 <= _zz_b_45;
    _zz_b_47 <= _zz_b_46;
    _zz_b_48 <= _zz_b_47;
    _zz_b_49 <= _zz__zz_5_port1;
    _zz_b_50 <= _zz_b_49;
    _zz_b_51 <= _zz_b_50;
    _zz_b_52 <= _zz_b_51;
    _zz_b_53 <= _zz_b_52;
    _zz_b_54 <= _zz_b_53;
    _zz_b_55 <= _zz_b_54;
    _zz_b_56 <= _zz_b_55;
    _zz_b_57 <= _zz_b_56;
    _zz_b_58 <= _zz_b_57;
    _zz_b_59 <= _zz__zz_6_port1;
    _zz_b_60 <= _zz_b_59;
    _zz_b_61 <= _zz_b_60;
    _zz_b_62 <= _zz_b_61;
    _zz_b_63 <= _zz_b_62;
    _zz_b_64 <= _zz_b_63;
    _zz_b_65 <= _zz_b_64;
    _zz_b_66 <= _zz_b_65;
    _zz_b_67 <= _zz_b_66;
    _zz_b_68 <= _zz_b_67;
    _zz_b_69 <= _zz__zz_7_port1;
    _zz_b_70 <= _zz_b_69;
    _zz_b_71 <= _zz_b_70;
    _zz_b_72 <= _zz_b_71;
    _zz_b_73 <= _zz_b_72;
    _zz_b_74 <= _zz_b_73;
    _zz_b_75 <= _zz_b_74;
    _zz_b_76 <= _zz_b_75;
    _zz_b_77 <= _zz_b_76;
    _zz_b_78 <= _zz_b_77;
    _zz_b_79 <= _zz__zz_8_port1;
    _zz_b_80 <= _zz_b_79;
    _zz_b_81 <= _zz_b_80;
    _zz_b_82 <= _zz_b_81;
    _zz_b_83 <= _zz_b_82;
    _zz_b_84 <= _zz_b_83;
    _zz_b_85 <= _zz_b_84;
    _zz_b_86 <= _zz_b_85;
    _zz_b_87 <= _zz_b_86;
    _zz_b_88 <= _zz_b_87;
    _zz_b_89 <= _zz__zz_9_port1;
    _zz_b_90 <= _zz_b_89;
    _zz_b_91 <= _zz_b_90;
    _zz_b_92 <= _zz_b_91;
    _zz_b_93 <= _zz_b_92;
    _zz_b_94 <= _zz_b_93;
    _zz_b_95 <= _zz_b_94;
    _zz_b_96 <= _zz_b_95;
    _zz_b_97 <= _zz_b_96;
    _zz_b_98 <= _zz_b_97;
  end


endmodule

module ConvState (
  input      [3:0]    control,
  input      [3:0]    complete,
  output reg [3:0]    state,
  output reg [3:0]    sign,
  output reg          dmaReadValid,
  output reg          dmaWriteValid,
  output reg          softReset,
  input               clk,
  input               reset
);
  localparam ConvStateEnum_IDLE = 5'd1;
  localparam ConvStateEnum_PARA = 5'd2;
  localparam ConvStateEnum_PARA_IRQ = 5'd4;
  localparam ConvStateEnum_COMPUTE = 5'd8;
  localparam ConvStateEnum_COMPUTE_IRQ = 5'd16;

  reg        [4:0]    fsm_currentState;
  reg        [4:0]    fsm_nextState;
  wire                when_ConvState_l80;
  wire                when_ConvState_l82;
  wire                when_ConvState_l89;
  wire                when_ConvState_l96;
  wire                when_ConvState_l103;
  wire                when_ConvState_l110;
  reg                 dmaReadValid_1;
  reg                 dmaWriteValid_1;
  reg                 dmaWriteValid_1_delay_1;
  reg                 dmaWriteValid_1_delay_2;
  reg                 dmaWriteValid_1_delay_3;
  reg                 dmaWriteValid_1_delay_4;
  reg                 dmaReadValid_1_delay_1;
  reg                 dmaReadValid_1_delay_2;
  reg                 dmaReadValid_1_delay_3;
  reg                 dmaReadValid_1_delay_4;
  wire                when_ConvState_l157;
  wire                when_ConvState_l161;
  wire                when_ConvState_l171;
  `ifndef SYNTHESIS
  reg [87:0] fsm_currentState_string;
  reg [87:0] fsm_nextState_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      ConvStateEnum_IDLE : fsm_currentState_string = "IDLE       ";
      ConvStateEnum_PARA : fsm_currentState_string = "PARA       ";
      ConvStateEnum_PARA_IRQ : fsm_currentState_string = "PARA_IRQ   ";
      ConvStateEnum_COMPUTE : fsm_currentState_string = "COMPUTE    ";
      ConvStateEnum_COMPUTE_IRQ : fsm_currentState_string = "COMPUTE_IRQ";
      default : fsm_currentState_string = "???????????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      ConvStateEnum_IDLE : fsm_nextState_string = "IDLE       ";
      ConvStateEnum_PARA : fsm_nextState_string = "PARA       ";
      ConvStateEnum_PARA_IRQ : fsm_nextState_string = "PARA_IRQ   ";
      ConvStateEnum_COMPUTE : fsm_nextState_string = "COMPUTE    ";
      ConvStateEnum_COMPUTE_IRQ : fsm_nextState_string = "COMPUTE_IRQ";
      default : fsm_nextState_string = "???????????";
    endcase
  end
  `endif

  assign when_ConvState_l80 = (control == 4'b0001);
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & ConvStateEnum_IDLE) == ConvStateEnum_IDLE) : begin
        if(when_ConvState_l80) begin
          fsm_nextState = ConvStateEnum_PARA;
        end else begin
          if(when_ConvState_l82) begin
            fsm_nextState = ConvStateEnum_COMPUTE;
          end else begin
            fsm_nextState = ConvStateEnum_IDLE;
          end
        end
      end
      (((fsm_currentState) & ConvStateEnum_PARA) == ConvStateEnum_PARA) : begin
        if(when_ConvState_l89) begin
          fsm_nextState = ConvStateEnum_PARA_IRQ;
        end else begin
          fsm_nextState = ConvStateEnum_PARA;
        end
      end
      (((fsm_currentState) & ConvStateEnum_PARA_IRQ) == ConvStateEnum_PARA_IRQ) : begin
        if(when_ConvState_l96) begin
          fsm_nextState = ConvStateEnum_IDLE;
        end else begin
          fsm_nextState = ConvStateEnum_PARA_IRQ;
        end
      end
      (((fsm_currentState) & ConvStateEnum_COMPUTE) == ConvStateEnum_COMPUTE) : begin
        if(when_ConvState_l103) begin
          fsm_nextState = ConvStateEnum_COMPUTE_IRQ;
        end else begin
          fsm_nextState = ConvStateEnum_COMPUTE;
        end
      end
      default : begin
        if(when_ConvState_l110) begin
          fsm_nextState = ConvStateEnum_IDLE;
        end else begin
          fsm_nextState = ConvStateEnum_COMPUTE_IRQ;
        end
      end
    endcase
  end

  assign when_ConvState_l82 = (control == 4'b0010);
  assign when_ConvState_l89 = (complete == 4'b0001);
  assign when_ConvState_l96 = (control == 4'b1111);
  assign when_ConvState_l103 = (complete == 4'b0010);
  assign when_ConvState_l110 = (control == 4'b1111);
  assign when_ConvState_l157 = (((fsm_currentState & ConvStateEnum_IDLE) != 5'b00000) && ((fsm_nextState & ConvStateEnum_PARA) != 5'b00000));
  assign when_ConvState_l161 = (((fsm_currentState & ConvStateEnum_IDLE) != 5'b00000) && ((fsm_nextState & ConvStateEnum_COMPUTE) != 5'b00000));
  assign when_ConvState_l171 = (((fsm_currentState & ConvStateEnum_COMPUTE_IRQ) != 5'b00000) && ((fsm_nextState & ConvStateEnum_IDLE) != 5'b00000));
  always @(*) begin
    if(when_ConvState_l171) begin
      softReset = 1'b1;
    end else begin
      softReset = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      dmaReadValid <= 1'b0;
      dmaWriteValid <= 1'b0;
      fsm_currentState <= ConvStateEnum_IDLE;
      dmaReadValid_1 <= 1'b0;
      dmaWriteValid_1 <= 1'b0;
    end else begin
      fsm_currentState <= fsm_nextState;
      dmaWriteValid <= dmaWriteValid_1_delay_4;
      dmaReadValid <= dmaReadValid_1_delay_4;
      if(when_ConvState_l157) begin
        dmaReadValid_1 <= 1'b1;
        dmaWriteValid_1 <= 1'b0;
      end else begin
        if(when_ConvState_l161) begin
          dmaWriteValid_1 <= 1'b1;
          dmaReadValid_1 <= 1'b1;
        end else begin
          dmaReadValid_1 <= 1'b0;
          dmaWriteValid_1 <= 1'b0;
        end
      end
    end
  end

  always @(posedge clk) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & ConvStateEnum_IDLE) == ConvStateEnum_IDLE) : begin
        state <= 4'b0000;
      end
      (((fsm_currentState) & ConvStateEnum_PARA) == ConvStateEnum_PARA) : begin
        state <= 4'b0001;
      end
      (((fsm_currentState) & ConvStateEnum_COMPUTE) == ConvStateEnum_COMPUTE) : begin
        state <= 4'b0010;
      end
      (((fsm_currentState) & ConvStateEnum_COMPUTE_IRQ) == ConvStateEnum_COMPUTE_IRQ) : begin
        state <= 4'b1111;
      end
      default : begin
        state <= 4'b1111;
      end
    endcase
    dmaWriteValid_1_delay_1 <= dmaWriteValid_1;
    dmaWriteValid_1_delay_2 <= dmaWriteValid_1_delay_1;
    dmaWriteValid_1_delay_3 <= dmaWriteValid_1_delay_2;
    dmaWriteValid_1_delay_4 <= dmaWriteValid_1_delay_3;
    dmaReadValid_1_delay_1 <= dmaReadValid_1;
    dmaReadValid_1_delay_2 <= dmaReadValid_1_delay_1;
    dmaReadValid_1_delay_3 <= dmaReadValid_1_delay_2;
    dmaReadValid_1_delay_4 <= dmaReadValid_1_delay_3;
    if(when_ConvState_l157) begin
      sign <= 4'b0001;
    end else begin
      if(when_ConvState_l161) begin
        sign <= 4'b0010;
      end else begin
        sign <= 4'b0000;
      end
    end
  end


endmodule

module Stride (
  input               sData_valid,
  output reg          sData_ready,
  input      [127:0]  sData_payload,
  output              mData_valid,
  input               mData_ready,
  output     [127:0]  mData_payload,
  output reg          sReady,
  output              complete,
  input               enStride,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input      [11:0]   channelOut,
  input               start,
  output              last,
  input               clk,
  input               reset,
  input               softReset
);
  localparam StrideEnum_IDLE = 3'd1;
  localparam StrideEnum_INIT = 3'd2;
  localparam StrideEnum_STRIDE = 3'd4;

  reg                 fifo_push_valid;
  wire                fifo_push_ready;
  wire                fifo_pop_valid;
  wire       [127:0]  fifo_pop_payload;
  wire       [14:0]   fifo_availability;
  wire       [7:0]    _zz_when_WaCounter_l12_1;
  wire       [9:0]    _zz_when_WaCounter_l12_2;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire       [17:0]   _zz_when_Stride_l99;
  wire       [8:0]    _zz_colOutTimes;
  wire       [8:0]    _zz_rowOutTimes;
  wire       [7:0]    _zz_when_WaCounter_l12_4;
  wire       [9:0]    _zz_when_WaCounter_l12_5;
  wire       [9:0]    _zz_when_WaCounter_l12_6;
  wire                fsm_initEnd;
  reg        [2:0]    fsm_currentState;
  reg        [2:0]    fsm_nextState;
  wire                when_WaCounter_l17;
  reg        [2:0]    initCnt_count;
  reg                 initCnt_valid;
  wire                when_WaCounter_l12;
  wire                when_Stride_l67;
  reg        [7:0]    channelTimes;
  wire                when_Stride_l68;
  reg        [9:0]    colTimes;
  wire                when_Stride_l69;
  reg        [9:0]    rowTimes;
  reg        [17:0]   dataCount;
  wire                sData_fire;
  wire                when_WaCounter_l17_1;
  reg        [7:0]    channelCnt_count;
  reg                 channelCnt_valid;
  wire                when_WaCounter_l12_1;
  wire                sData_fire_1;
  wire                when_WaCounter_l17_2;
  reg        [9:0]    colCnt_count;
  reg                 colCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                sData_fire_2;
  wire                when_WaCounter_l17_3;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                sData_fire_3;
  wire                when_Stride_l80;
  wire                when_Stride_l86;
  wire                when_Stream_l438;
  reg                 sData_thrown_valid;
  wire                sData_thrown_ready;
  wire                when_Stride_l99;
  reg        [9:0]    colOutTimes;
  reg        [9:0]    rowOutTimes;
  wire                mData_fire;
  reg        [7:0]    channelOutCnt_count;
  reg                 channelOutCnt_valid;
  wire                when_WaCounter_l12_4;
  wire                mData_fire_1;
  wire                when_WaCounter_l17_4;
  reg        [9:0]    colOutCnt_count;
  reg                 colOutCnt_valid;
  wire                when_WaCounter_l12_5;
  wire                mData_fire_2;
  wire                when_WaCounter_l17_5;
  reg        [9:0]    rowOutCnt_count;
  reg                 rowOutCnt_valid;
  wire                when_WaCounter_l12_6;
  `ifndef SYNTHESIS
  reg [47:0] fsm_currentState_string;
  reg [47:0] fsm_nextState_string;
  `endif


  assign _zz_when_WaCounter_l12_1 = (channelTimes - 8'h01);
  assign _zz_when_WaCounter_l12_2 = (colTimes - 10'h001);
  assign _zz_when_WaCounter_l12_3 = (rowTimes - 10'h001);
  assign _zz_when_Stride_l99 = {3'd0, fifo_availability};
  assign _zz_colOutTimes = (colTimes >>> 1);
  assign _zz_rowOutTimes = (rowTimes >>> 1);
  assign _zz_when_WaCounter_l12_4 = (channelTimes - 8'h01);
  assign _zz_when_WaCounter_l12_5 = (colOutTimes - 10'h001);
  assign _zz_when_WaCounter_l12_6 = (rowOutTimes - 10'h001);
  WaStreamFifoPipe fifo (
    .push_valid   (fifo_push_valid        ), //i
    .push_ready   (fifo_push_ready        ), //o
    .push_payload (sData_payload[127:0]   ), //i
    .pop_valid    (fifo_pop_valid         ), //o
    .pop_ready    (mData_ready            ), //i
    .pop_payload  (fifo_pop_payload[127:0]), //o
    .flush        (1'b0                   ), //i
    .availability (fifo_availability[14:0]), //o
    .clk          (clk                    ), //i
    .reset        (reset                  ), //i
    .softReset    (softReset              )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      StrideEnum_IDLE : fsm_currentState_string = "IDLE  ";
      StrideEnum_INIT : fsm_currentState_string = "INIT  ";
      StrideEnum_STRIDE : fsm_currentState_string = "STRIDE";
      default : fsm_currentState_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      StrideEnum_IDLE : fsm_nextState_string = "IDLE  ";
      StrideEnum_INIT : fsm_nextState_string = "INIT  ";
      StrideEnum_STRIDE : fsm_nextState_string = "STRIDE";
      default : fsm_nextState_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & StrideEnum_IDLE) == StrideEnum_IDLE) : begin
        if(start) begin
          fsm_nextState = StrideEnum_INIT;
        end else begin
          fsm_nextState = StrideEnum_IDLE;
        end
      end
      (((fsm_currentState) & StrideEnum_INIT) == StrideEnum_INIT) : begin
        if(fsm_initEnd) begin
          fsm_nextState = StrideEnum_STRIDE;
        end else begin
          fsm_nextState = StrideEnum_INIT;
        end
      end
      default : begin
        if(complete) begin
          fsm_nextState = StrideEnum_IDLE;
        end else begin
          fsm_nextState = StrideEnum_STRIDE;
        end
      end
    endcase
  end

  assign when_WaCounter_l17 = ((fsm_currentState & StrideEnum_INIT) != 3'b000);
  assign when_WaCounter_l12 = (initCnt_count == 3'b111);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCnt_valid = 1'b1;
    end else begin
      initCnt_valid = 1'b0;
    end
    if(when_Stride_l80) begin
      initCnt_valid = 1'b0;
    end
  end

  assign fsm_initEnd = initCnt_valid;
  assign when_Stride_l67 = ((fsm_currentState & StrideEnum_INIT) != 3'b000);
  assign when_Stride_l68 = ((fsm_currentState & StrideEnum_INIT) != 3'b000);
  assign when_Stride_l69 = ((fsm_currentState & StrideEnum_INIT) != 3'b000);
  assign sData_fire = (sData_valid && sData_ready);
  assign when_WaCounter_l17_1 = (((fsm_currentState & StrideEnum_STRIDE) != 3'b000) && sData_fire);
  assign when_WaCounter_l12_1 = (channelCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelCnt_valid = 1'b1;
    end else begin
      channelCnt_valid = 1'b0;
    end
    if(when_Stride_l80) begin
      channelCnt_valid = 1'b0;
    end
  end

  assign sData_fire_1 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_2 = (channelCnt_valid && sData_fire_1);
  assign when_WaCounter_l12_2 = (colCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      colCnt_valid = 1'b1;
    end else begin
      colCnt_valid = 1'b0;
    end
    if(when_Stride_l80) begin
      colCnt_valid = 1'b0;
    end
  end

  assign sData_fire_2 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_3 = ((channelCnt_valid && colCnt_valid) && sData_fire_2);
  assign when_WaCounter_l12_3 = (rowCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
    if(when_Stride_l80) begin
      rowCnt_valid = 1'b0;
    end
  end

  assign sData_fire_3 = (sData_valid && sData_ready);
  assign complete = (((rowCnt_valid && colCnt_valid) && channelCnt_valid) && sData_fire_3);
  assign when_Stride_l80 = ((fsm_currentState & StrideEnum_IDLE) != 3'b000);
  assign when_Stride_l86 = ((fsm_currentState & StrideEnum_STRIDE) != 3'b000);
  assign when_Stream_l438 = (colCnt_count[0] || rowCnt_count[0]);
  always @(*) begin
    sData_thrown_valid = sData_valid;
    if(when_Stream_l438) begin
      sData_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_Stride_l86) begin
      if(enStride) begin
        sData_ready = sData_thrown_ready;
        if(when_Stream_l438) begin
          sData_ready = 1'b1;
        end
      end else begin
        sData_ready = fifo_push_ready;
      end
    end else begin
      sData_ready = 1'b0;
    end
  end

  always @(*) begin
    if(when_Stride_l86) begin
      if(enStride) begin
        fifo_push_valid = sData_thrown_valid;
      end else begin
        fifo_push_valid = sData_valid;
      end
    end else begin
      fifo_push_valid = 1'b0;
    end
  end

  assign sData_thrown_ready = fifo_push_ready;
  assign when_Stride_l99 = (dataCount < _zz_when_Stride_l99);
  always @(*) begin
    if(when_Stride_l99) begin
      sReady = 1'b1;
    end else begin
      sReady = 1'b0;
    end
  end

  assign mData_valid = fifo_pop_valid;
  assign mData_payload = fifo_pop_payload;
  assign mData_fire = (mData_valid && mData_ready);
  assign when_WaCounter_l12_4 = (channelOutCnt_count == _zz_when_WaCounter_l12_4);
  always @(*) begin
    if(when_WaCounter_l12_4) begin
      channelOutCnt_valid = 1'b1;
    end else begin
      channelOutCnt_valid = 1'b0;
    end
  end

  assign mData_fire_1 = (mData_valid && mData_ready);
  assign when_WaCounter_l17_4 = (channelOutCnt_valid && mData_fire_1);
  assign when_WaCounter_l12_5 = (colOutCnt_count == _zz_when_WaCounter_l12_5);
  always @(*) begin
    if(when_WaCounter_l12_5) begin
      colOutCnt_valid = 1'b1;
    end else begin
      colOutCnt_valid = 1'b0;
    end
  end

  assign mData_fire_2 = (mData_valid && mData_ready);
  assign when_WaCounter_l17_5 = ((channelOutCnt_valid && colOutCnt_valid) && mData_fire_2);
  assign when_WaCounter_l12_6 = (rowOutCnt_count == _zz_when_WaCounter_l12_6);
  always @(*) begin
    if(when_WaCounter_l12_6) begin
      rowOutCnt_valid = 1'b1;
    end else begin
      rowOutCnt_valid = 1'b0;
    end
  end

  assign last = ((channelOutCnt_valid && colOutCnt_valid) && rowOutCnt_valid);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      fsm_currentState <= StrideEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 8'h0;
      colCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      channelOutCnt_count <= 8'h0;
      colOutCnt_count <= 10'h0;
      rowOutCnt_count <= 10'h0;
    end else begin
      if(softReset) begin
      fsm_currentState <= StrideEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 8'h0;
      colCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      channelOutCnt_count <= 8'h0;
      colOutCnt_count <= 10'h0;
      rowOutCnt_count <= 10'h0;
      end else begin
        fsm_currentState <= fsm_nextState;
        if(when_WaCounter_l17) begin
          initCnt_count <= (initCnt_count + 3'b001);
          if(initCnt_valid) begin
            initCnt_count <= 3'b000;
          end
        end
        if(when_WaCounter_l17_1) begin
          channelCnt_count <= (channelCnt_count + 8'h01);
          if(channelCnt_valid) begin
            channelCnt_count <= 8'h0;
          end
        end
        if(when_WaCounter_l17_2) begin
          colCnt_count <= (colCnt_count + 10'h001);
          if(colCnt_valid) begin
            colCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_3) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
        if(when_Stride_l80) begin
          initCnt_count <= 3'b000;
          channelCnt_count <= 8'h0;
          colCnt_count <= 10'h0;
          rowCnt_count <= 10'h0;
        end
        if(mData_fire) begin
          channelOutCnt_count <= (channelOutCnt_count + 8'h01);
          if(channelOutCnt_valid) begin
            channelOutCnt_count <= 8'h0;
          end
        end
        if(when_WaCounter_l17_4) begin
          colOutCnt_count <= (colOutCnt_count + 10'h001);
          if(colOutCnt_valid) begin
            colOutCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_5) begin
          rowOutCnt_count <= (rowOutCnt_count + 10'h001);
          if(rowOutCnt_valid) begin
            rowOutCnt_count <= 10'h0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(when_Stride_l67) begin
      channelTimes <= (channelOut >>> 4);
    end
    if(when_Stride_l68) begin
      colTimes <= colNumIn;
    end
    if(when_Stride_l69) begin
      rowTimes <= rowNumIn;
    end
    dataCount <= (channelTimes * colTimes);
    if(enStride) begin
      colOutTimes <= {1'd0, _zz_colOutTimes};
      rowOutTimes <= {1'd0, _zz_rowOutTimes};
    end else begin
      colOutTimes <= colTimes;
      rowOutTimes <= rowTimes;
    end
  end


endmodule

module Quan (
  input      [31:0]   dataIn_0,
  input      [31:0]   dataIn_1,
  input      [31:0]   dataIn_2,
  input      [31:0]   dataIn_3,
  input      [31:0]   dataIn_4,
  input      [31:0]   dataIn_5,
  input      [31:0]   dataIn_6,
  input      [31:0]   dataIn_7,
  input      [31:0]   dataIn_8,
  input      [31:0]   dataIn_9,
  input      [31:0]   dataIn_10,
  input      [31:0]   dataIn_11,
  input      [31:0]   dataIn_12,
  input      [31:0]   dataIn_13,
  input      [31:0]   dataIn_14,
  input      [31:0]   dataIn_15,
  input      [511:0]  biasIn,
  input      [511:0]  scaleIn,
  input      [511:0]  shiftIn,
  input      [7:0]    zeroIn,
  input               activationEn,
  output reg [127:0]  dataOut,
  input      [31:0]   amendReg,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [31:0]   bias_1_Bias_quan_0;
  wire       [31:0]   bias_1_Bias_quan_1;
  wire       [31:0]   bias_1_Bias_quan_2;
  wire       [31:0]   bias_1_Bias_quan_3;
  wire       [31:0]   bias_1_Bias_quan_4;
  wire       [31:0]   bias_1_Bias_quan_5;
  wire       [31:0]   bias_1_Bias_quan_6;
  wire       [31:0]   bias_1_Bias_quan_7;
  wire       [31:0]   bias_1_Bias_quan_8;
  wire       [31:0]   bias_1_Bias_quan_9;
  wire       [31:0]   bias_1_Bias_quan_10;
  wire       [31:0]   bias_1_Bias_quan_11;
  wire       [31:0]   bias_1_Bias_quan_12;
  wire       [31:0]   bias_1_Bias_quan_13;
  wire       [31:0]   bias_1_Bias_quan_14;
  wire       [31:0]   bias_1_Bias_quan_15;
  wire       [47:0]   bias_1_Bias_dataOut_0;
  wire       [47:0]   bias_1_Bias_dataOut_1;
  wire       [47:0]   bias_1_Bias_dataOut_2;
  wire       [47:0]   bias_1_Bias_dataOut_3;
  wire       [47:0]   bias_1_Bias_dataOut_4;
  wire       [47:0]   bias_1_Bias_dataOut_5;
  wire       [47:0]   bias_1_Bias_dataOut_6;
  wire       [47:0]   bias_1_Bias_dataOut_7;
  wire       [47:0]   bias_1_Bias_dataOut_8;
  wire       [47:0]   bias_1_Bias_dataOut_9;
  wire       [47:0]   bias_1_Bias_dataOut_10;
  wire       [47:0]   bias_1_Bias_dataOut_11;
  wire       [47:0]   bias_1_Bias_dataOut_12;
  wire       [47:0]   bias_1_Bias_dataOut_13;
  wire       [47:0]   bias_1_Bias_dataOut_14;
  wire       [47:0]   bias_1_Bias_dataOut_15;
  wire       [31:0]   scale_1_Scale_dataOut_0;
  wire       [31:0]   scale_1_Scale_dataOut_1;
  wire       [31:0]   scale_1_Scale_dataOut_2;
  wire       [31:0]   scale_1_Scale_dataOut_3;
  wire       [31:0]   scale_1_Scale_dataOut_4;
  wire       [31:0]   scale_1_Scale_dataOut_5;
  wire       [31:0]   scale_1_Scale_dataOut_6;
  wire       [31:0]   scale_1_Scale_dataOut_7;
  wire       [31:0]   scale_1_Scale_dataOut_8;
  wire       [31:0]   scale_1_Scale_dataOut_9;
  wire       [31:0]   scale_1_Scale_dataOut_10;
  wire       [31:0]   scale_1_Scale_dataOut_11;
  wire       [31:0]   scale_1_Scale_dataOut_12;
  wire       [31:0]   scale_1_Scale_dataOut_13;
  wire       [31:0]   scale_1_Scale_dataOut_14;
  wire       [31:0]   scale_1_Scale_dataOut_15;
  wire       [15:0]   shift_1_shift_dataOut_0;
  wire       [15:0]   shift_1_shift_dataOut_1;
  wire       [15:0]   shift_1_shift_dataOut_2;
  wire       [15:0]   shift_1_shift_dataOut_3;
  wire       [15:0]   shift_1_shift_dataOut_4;
  wire       [15:0]   shift_1_shift_dataOut_5;
  wire       [15:0]   shift_1_shift_dataOut_6;
  wire       [15:0]   shift_1_shift_dataOut_7;
  wire       [15:0]   shift_1_shift_dataOut_8;
  wire       [15:0]   shift_1_shift_dataOut_9;
  wire       [15:0]   shift_1_shift_dataOut_10;
  wire       [15:0]   shift_1_shift_dataOut_11;
  wire       [15:0]   shift_1_shift_dataOut_12;
  wire       [15:0]   shift_1_shift_dataOut_13;
  wire       [15:0]   shift_1_shift_dataOut_14;
  wire       [15:0]   shift_1_shift_dataOut_15;
  wire       [7:0]    zero_1_dataOut_0;
  wire       [7:0]    zero_1_dataOut_1;
  wire       [7:0]    zero_1_dataOut_2;
  wire       [7:0]    zero_1_dataOut_3;
  wire       [7:0]    zero_1_dataOut_4;
  wire       [7:0]    zero_1_dataOut_5;
  wire       [7:0]    zero_1_dataOut_6;
  wire       [7:0]    zero_1_dataOut_7;
  wire       [7:0]    zero_1_dataOut_8;
  wire       [7:0]    zero_1_dataOut_9;
  wire       [7:0]    zero_1_dataOut_10;
  wire       [7:0]    zero_1_dataOut_11;
  wire       [7:0]    zero_1_dataOut_12;
  wire       [7:0]    zero_1_dataOut_13;
  wire       [7:0]    zero_1_dataOut_14;
  wire       [7:0]    zero_1_dataOut_15;
  wire       [7:0]    leakyRelu_1_dataOut_0;
  wire       [7:0]    leakyRelu_1_dataOut_1;
  wire       [7:0]    leakyRelu_1_dataOut_2;
  wire       [7:0]    leakyRelu_1_dataOut_3;
  wire       [7:0]    leakyRelu_1_dataOut_4;
  wire       [7:0]    leakyRelu_1_dataOut_5;
  wire       [7:0]    leakyRelu_1_dataOut_6;
  wire       [7:0]    leakyRelu_1_dataOut_7;
  wire       [7:0]    leakyRelu_1_dataOut_8;
  wire       [7:0]    leakyRelu_1_dataOut_9;
  wire       [7:0]    leakyRelu_1_dataOut_10;
  wire       [7:0]    leakyRelu_1_dataOut_11;
  wire       [7:0]    leakyRelu_1_dataOut_12;
  wire       [7:0]    leakyRelu_1_dataOut_13;
  wire       [7:0]    leakyRelu_1_dataOut_14;
  wire       [7:0]    leakyRelu_1_dataOut_15;
  reg        [31:0]   dataIn_regNext_0;
  reg        [31:0]   dataIn_regNext_1;
  reg        [31:0]   dataIn_regNext_2;
  reg        [31:0]   dataIn_regNext_3;
  reg        [31:0]   dataIn_regNext_4;
  reg        [31:0]   dataIn_regNext_5;
  reg        [31:0]   dataIn_regNext_6;
  reg        [31:0]   dataIn_regNext_7;
  reg        [31:0]   dataIn_regNext_8;
  reg        [31:0]   dataIn_regNext_9;
  reg        [31:0]   dataIn_regNext_10;
  reg        [31:0]   dataIn_regNext_11;
  reg        [31:0]   dataIn_regNext_12;
  reg        [31:0]   dataIn_regNext_13;
  reg        [31:0]   dataIn_regNext_14;
  reg        [31:0]   dataIn_regNext_15;
  reg        [31:0]   _zz_Scale_quan_0;
  reg        [31:0]   _zz_Scale_quan_1;
  reg        [31:0]   _zz_Scale_quan_2;
  reg        [31:0]   _zz_Scale_quan_3;
  reg        [31:0]   _zz_Scale_quan_4;
  reg        [31:0]   _zz_Scale_quan_5;
  reg        [31:0]   _zz_Scale_quan_6;
  reg        [31:0]   _zz_Scale_quan_7;
  reg        [31:0]   _zz_Scale_quan_8;
  reg        [31:0]   _zz_Scale_quan_9;
  reg        [31:0]   _zz_Scale_quan_10;
  reg        [31:0]   _zz_Scale_quan_11;
  reg        [31:0]   _zz_Scale_quan_12;
  reg        [31:0]   _zz_Scale_quan_13;
  reg        [31:0]   _zz_Scale_quan_14;
  reg        [31:0]   _zz_Scale_quan_15;
  reg        [31:0]   _zz_Scale_quan_0_1;
  reg        [31:0]   _zz_Scale_quan_1_1;
  reg        [31:0]   _zz_Scale_quan_2_1;
  reg        [31:0]   _zz_Scale_quan_3_1;
  reg        [31:0]   _zz_Scale_quan_4_1;
  reg        [31:0]   _zz_Scale_quan_5_1;
  reg        [31:0]   _zz_Scale_quan_6_1;
  reg        [31:0]   _zz_Scale_quan_7_1;
  reg        [31:0]   _zz_Scale_quan_8_1;
  reg        [31:0]   _zz_Scale_quan_9_1;
  reg        [31:0]   _zz_Scale_quan_10_1;
  reg        [31:0]   _zz_Scale_quan_11_1;
  reg        [31:0]   _zz_Scale_quan_12_1;
  reg        [31:0]   _zz_Scale_quan_13_1;
  reg        [31:0]   _zz_Scale_quan_14_1;
  reg        [31:0]   _zz_Scale_quan_15_1;
  reg        [31:0]   _zz_shift_quan_0;
  reg        [31:0]   _zz_shift_quan_1;
  reg        [31:0]   _zz_shift_quan_2;
  reg        [31:0]   _zz_shift_quan_3;
  reg        [31:0]   _zz_shift_quan_4;
  reg        [31:0]   _zz_shift_quan_5;
  reg        [31:0]   _zz_shift_quan_6;
  reg        [31:0]   _zz_shift_quan_7;
  reg        [31:0]   _zz_shift_quan_8;
  reg        [31:0]   _zz_shift_quan_9;
  reg        [31:0]   _zz_shift_quan_10;
  reg        [31:0]   _zz_shift_quan_11;
  reg        [31:0]   _zz_shift_quan_12;
  reg        [31:0]   _zz_shift_quan_13;
  reg        [31:0]   _zz_shift_quan_14;
  reg        [31:0]   _zz_shift_quan_15;
  reg        [31:0]   _zz_shift_quan_0_1;
  reg        [31:0]   _zz_shift_quan_1_1;
  reg        [31:0]   _zz_shift_quan_2_1;
  reg        [31:0]   _zz_shift_quan_3_1;
  reg        [31:0]   _zz_shift_quan_4_1;
  reg        [31:0]   _zz_shift_quan_5_1;
  reg        [31:0]   _zz_shift_quan_6_1;
  reg        [31:0]   _zz_shift_quan_7_1;
  reg        [31:0]   _zz_shift_quan_8_1;
  reg        [31:0]   _zz_shift_quan_9_1;
  reg        [31:0]   _zz_shift_quan_10_1;
  reg        [31:0]   _zz_shift_quan_11_1;
  reg        [31:0]   _zz_shift_quan_12_1;
  reg        [31:0]   _zz_shift_quan_13_1;
  reg        [31:0]   _zz_shift_quan_14_1;
  reg        [31:0]   _zz_shift_quan_15_1;
  reg        [31:0]   _zz_shift_quan_0_2;
  reg        [31:0]   _zz_shift_quan_1_2;
  reg        [31:0]   _zz_shift_quan_2_2;
  reg        [31:0]   _zz_shift_quan_3_2;
  reg        [31:0]   _zz_shift_quan_4_2;
  reg        [31:0]   _zz_shift_quan_5_2;
  reg        [31:0]   _zz_shift_quan_6_2;
  reg        [31:0]   _zz_shift_quan_7_2;
  reg        [31:0]   _zz_shift_quan_8_2;
  reg        [31:0]   _zz_shift_quan_9_2;
  reg        [31:0]   _zz_shift_quan_10_2;
  reg        [31:0]   _zz_shift_quan_11_2;
  reg        [31:0]   _zz_shift_quan_12_2;
  reg        [31:0]   _zz_shift_quan_13_2;
  reg        [31:0]   _zz_shift_quan_14_2;
  reg        [31:0]   _zz_shift_quan_15_2;
  reg        [31:0]   _zz_shift_quan_0_3;
  reg        [31:0]   _zz_shift_quan_1_3;
  reg        [31:0]   _zz_shift_quan_2_3;
  reg        [31:0]   _zz_shift_quan_3_3;
  reg        [31:0]   _zz_shift_quan_4_3;
  reg        [31:0]   _zz_shift_quan_5_3;
  reg        [31:0]   _zz_shift_quan_6_3;
  reg        [31:0]   _zz_shift_quan_7_3;
  reg        [31:0]   _zz_shift_quan_8_3;
  reg        [31:0]   _zz_shift_quan_9_3;
  reg        [31:0]   _zz_shift_quan_10_3;
  reg        [31:0]   _zz_shift_quan_11_3;
  reg        [31:0]   _zz_shift_quan_12_3;
  reg        [31:0]   _zz_shift_quan_13_3;
  reg        [31:0]   _zz_shift_quan_14_3;
  reg        [31:0]   _zz_shift_quan_15_3;
  reg        [31:0]   _zz_shift_quan_0_4;
  reg        [31:0]   _zz_shift_quan_1_4;
  reg        [31:0]   _zz_shift_quan_2_4;
  reg        [31:0]   _zz_shift_quan_3_4;
  reg        [31:0]   _zz_shift_quan_4_4;
  reg        [31:0]   _zz_shift_quan_5_4;
  reg        [31:0]   _zz_shift_quan_6_4;
  reg        [31:0]   _zz_shift_quan_7_4;
  reg        [31:0]   _zz_shift_quan_8_4;
  reg        [31:0]   _zz_shift_quan_9_4;
  reg        [31:0]   _zz_shift_quan_10_4;
  reg        [31:0]   _zz_shift_quan_11_4;
  reg        [31:0]   _zz_shift_quan_12_4;
  reg        [31:0]   _zz_shift_quan_13_4;
  reg        [31:0]   _zz_shift_quan_14_4;
  reg        [31:0]   _zz_shift_quan_15_4;
  reg        [31:0]   _zz_shift_quan_0_5;
  reg        [31:0]   _zz_shift_quan_1_5;
  reg        [31:0]   _zz_shift_quan_2_5;
  reg        [31:0]   _zz_shift_quan_3_5;
  reg        [31:0]   _zz_shift_quan_4_5;
  reg        [31:0]   _zz_shift_quan_5_5;
  reg        [31:0]   _zz_shift_quan_6_5;
  reg        [31:0]   _zz_shift_quan_7_5;
  reg        [31:0]   _zz_shift_quan_8_5;
  reg        [31:0]   _zz_shift_quan_9_5;
  reg        [31:0]   _zz_shift_quan_10_5;
  reg        [31:0]   _zz_shift_quan_11_5;
  reg        [31:0]   _zz_shift_quan_12_5;
  reg        [31:0]   _zz_shift_quan_13_5;
  reg        [31:0]   _zz_shift_quan_14_5;
  reg        [31:0]   _zz_shift_quan_15_5;
  reg        [31:0]   _zz_shift_quan_0_6;
  reg        [31:0]   _zz_shift_quan_1_6;
  reg        [31:0]   _zz_shift_quan_2_6;
  reg        [31:0]   _zz_shift_quan_3_6;
  reg        [31:0]   _zz_shift_quan_4_6;
  reg        [31:0]   _zz_shift_quan_5_6;
  reg        [31:0]   _zz_shift_quan_6_6;
  reg        [31:0]   _zz_shift_quan_7_6;
  reg        [31:0]   _zz_shift_quan_8_6;
  reg        [31:0]   _zz_shift_quan_9_6;
  reg        [31:0]   _zz_shift_quan_10_6;
  reg        [31:0]   _zz_shift_quan_11_6;
  reg        [31:0]   _zz_shift_quan_12_6;
  reg        [31:0]   _zz_shift_quan_13_6;
  reg        [31:0]   _zz_shift_quan_14_6;
  reg        [31:0]   _zz_shift_quan_15_6;
  reg        [31:0]   _zz_shift_quan_0_7;
  reg        [31:0]   _zz_shift_quan_1_7;
  reg        [31:0]   _zz_shift_quan_2_7;
  reg        [31:0]   _zz_shift_quan_3_7;
  reg        [31:0]   _zz_shift_quan_4_7;
  reg        [31:0]   _zz_shift_quan_5_7;
  reg        [31:0]   _zz_shift_quan_6_7;
  reg        [31:0]   _zz_shift_quan_7_7;
  reg        [31:0]   _zz_shift_quan_8_7;
  reg        [31:0]   _zz_shift_quan_9_7;
  reg        [31:0]   _zz_shift_quan_10_7;
  reg        [31:0]   _zz_shift_quan_11_7;
  reg        [31:0]   _zz_shift_quan_12_7;
  reg        [31:0]   _zz_shift_quan_13_7;
  reg        [31:0]   _zz_shift_quan_14_7;
  reg        [31:0]   _zz_shift_quan_15_7;
  reg        [31:0]   _zz_shift_quan_0_8;
  reg        [31:0]   _zz_shift_quan_1_8;
  reg        [31:0]   _zz_shift_quan_2_8;
  reg        [31:0]   _zz_shift_quan_3_8;
  reg        [31:0]   _zz_shift_quan_4_8;
  reg        [31:0]   _zz_shift_quan_5_8;
  reg        [31:0]   _zz_shift_quan_6_8;
  reg        [31:0]   _zz_shift_quan_7_8;
  reg        [31:0]   _zz_shift_quan_8_8;
  reg        [31:0]   _zz_shift_quan_9_8;
  reg        [31:0]   _zz_shift_quan_10_8;
  reg        [31:0]   _zz_shift_quan_11_8;
  reg        [31:0]   _zz_shift_quan_12_8;
  reg        [31:0]   _zz_shift_quan_13_8;
  reg        [31:0]   _zz_shift_quan_14_8;
  reg        [31:0]   _zz_shift_quan_15_8;
  reg        [31:0]   _zz_shift_quan_0_9;
  reg        [31:0]   _zz_shift_quan_1_9;
  reg        [31:0]   _zz_shift_quan_2_9;
  reg        [31:0]   _zz_shift_quan_3_9;
  reg        [31:0]   _zz_shift_quan_4_9;
  reg        [31:0]   _zz_shift_quan_5_9;
  reg        [31:0]   _zz_shift_quan_6_9;
  reg        [31:0]   _zz_shift_quan_7_9;
  reg        [31:0]   _zz_shift_quan_8_9;
  reg        [31:0]   _zz_shift_quan_9_9;
  reg        [31:0]   _zz_shift_quan_10_9;
  reg        [31:0]   _zz_shift_quan_11_9;
  reg        [31:0]   _zz_shift_quan_12_9;
  reg        [31:0]   _zz_shift_quan_13_9;
  reg        [31:0]   _zz_shift_quan_14_9;
  reg        [31:0]   _zz_shift_quan_15_9;
  reg        [31:0]   _zz_shift_quan_0_10;
  reg        [31:0]   _zz_shift_quan_1_10;
  reg        [31:0]   _zz_shift_quan_2_10;
  reg        [31:0]   _zz_shift_quan_3_10;
  reg        [31:0]   _zz_shift_quan_4_10;
  reg        [31:0]   _zz_shift_quan_5_10;
  reg        [31:0]   _zz_shift_quan_6_10;
  reg        [31:0]   _zz_shift_quan_7_10;
  reg        [31:0]   _zz_shift_quan_8_10;
  reg        [31:0]   _zz_shift_quan_9_10;
  reg        [31:0]   _zz_shift_quan_10_10;
  reg        [31:0]   _zz_shift_quan_11_10;
  reg        [31:0]   _zz_shift_quan_12_10;
  reg        [31:0]   _zz_shift_quan_13_10;
  reg        [31:0]   _zz_shift_quan_14_10;
  reg        [31:0]   _zz_shift_quan_15_10;

  Bias bias_1 (
    .Bias_dataIn_0   (dataIn_regNext_0[31:0]      ), //i
    .Bias_dataIn_1   (dataIn_regNext_1[31:0]      ), //i
    .Bias_dataIn_2   (dataIn_regNext_2[31:0]      ), //i
    .Bias_dataIn_3   (dataIn_regNext_3[31:0]      ), //i
    .Bias_dataIn_4   (dataIn_regNext_4[31:0]      ), //i
    .Bias_dataIn_5   (dataIn_regNext_5[31:0]      ), //i
    .Bias_dataIn_6   (dataIn_regNext_6[31:0]      ), //i
    .Bias_dataIn_7   (dataIn_regNext_7[31:0]      ), //i
    .Bias_dataIn_8   (dataIn_regNext_8[31:0]      ), //i
    .Bias_dataIn_9   (dataIn_regNext_9[31:0]      ), //i
    .Bias_dataIn_10  (dataIn_regNext_10[31:0]     ), //i
    .Bias_dataIn_11  (dataIn_regNext_11[31:0]     ), //i
    .Bias_dataIn_12  (dataIn_regNext_12[31:0]     ), //i
    .Bias_dataIn_13  (dataIn_regNext_13[31:0]     ), //i
    .Bias_dataIn_14  (dataIn_regNext_14[31:0]     ), //i
    .Bias_dataIn_15  (dataIn_regNext_15[31:0]     ), //i
    .Bias_quan_0     (bias_1_Bias_quan_0[31:0]    ), //i
    .Bias_quan_1     (bias_1_Bias_quan_1[31:0]    ), //i
    .Bias_quan_2     (bias_1_Bias_quan_2[31:0]    ), //i
    .Bias_quan_3     (bias_1_Bias_quan_3[31:0]    ), //i
    .Bias_quan_4     (bias_1_Bias_quan_4[31:0]    ), //i
    .Bias_quan_5     (bias_1_Bias_quan_5[31:0]    ), //i
    .Bias_quan_6     (bias_1_Bias_quan_6[31:0]    ), //i
    .Bias_quan_7     (bias_1_Bias_quan_7[31:0]    ), //i
    .Bias_quan_8     (bias_1_Bias_quan_8[31:0]    ), //i
    .Bias_quan_9     (bias_1_Bias_quan_9[31:0]    ), //i
    .Bias_quan_10    (bias_1_Bias_quan_10[31:0]   ), //i
    .Bias_quan_11    (bias_1_Bias_quan_11[31:0]   ), //i
    .Bias_quan_12    (bias_1_Bias_quan_12[31:0]   ), //i
    .Bias_quan_13    (bias_1_Bias_quan_13[31:0]   ), //i
    .Bias_quan_14    (bias_1_Bias_quan_14[31:0]   ), //i
    .Bias_quan_15    (bias_1_Bias_quan_15[31:0]   ), //i
    .Bias_dataOut_0  (bias_1_Bias_dataOut_0[47:0] ), //o
    .Bias_dataOut_1  (bias_1_Bias_dataOut_1[47:0] ), //o
    .Bias_dataOut_2  (bias_1_Bias_dataOut_2[47:0] ), //o
    .Bias_dataOut_3  (bias_1_Bias_dataOut_3[47:0] ), //o
    .Bias_dataOut_4  (bias_1_Bias_dataOut_4[47:0] ), //o
    .Bias_dataOut_5  (bias_1_Bias_dataOut_5[47:0] ), //o
    .Bias_dataOut_6  (bias_1_Bias_dataOut_6[47:0] ), //o
    .Bias_dataOut_7  (bias_1_Bias_dataOut_7[47:0] ), //o
    .Bias_dataOut_8  (bias_1_Bias_dataOut_8[47:0] ), //o
    .Bias_dataOut_9  (bias_1_Bias_dataOut_9[47:0] ), //o
    .Bias_dataOut_10 (bias_1_Bias_dataOut_10[47:0]), //o
    .Bias_dataOut_11 (bias_1_Bias_dataOut_11[47:0]), //o
    .Bias_dataOut_12 (bias_1_Bias_dataOut_12[47:0]), //o
    .Bias_dataOut_13 (bias_1_Bias_dataOut_13[47:0]), //o
    .Bias_dataOut_14 (bias_1_Bias_dataOut_14[47:0]), //o
    .Bias_dataOut_15 (bias_1_Bias_dataOut_15[47:0]), //o
    .clk             (clk                         ), //i
    .reset           (reset                       ), //i
    .softReset       (softReset                   )  //i
  );
  Scale scale_1 (
    .Scale_dataIn_0   (bias_1_Bias_dataOut_0[47:0]   ), //i
    .Scale_dataIn_1   (bias_1_Bias_dataOut_1[47:0]   ), //i
    .Scale_dataIn_2   (bias_1_Bias_dataOut_2[47:0]   ), //i
    .Scale_dataIn_3   (bias_1_Bias_dataOut_3[47:0]   ), //i
    .Scale_dataIn_4   (bias_1_Bias_dataOut_4[47:0]   ), //i
    .Scale_dataIn_5   (bias_1_Bias_dataOut_5[47:0]   ), //i
    .Scale_dataIn_6   (bias_1_Bias_dataOut_6[47:0]   ), //i
    .Scale_dataIn_7   (bias_1_Bias_dataOut_7[47:0]   ), //i
    .Scale_dataIn_8   (bias_1_Bias_dataOut_8[47:0]   ), //i
    .Scale_dataIn_9   (bias_1_Bias_dataOut_9[47:0]   ), //i
    .Scale_dataIn_10  (bias_1_Bias_dataOut_10[47:0]  ), //i
    .Scale_dataIn_11  (bias_1_Bias_dataOut_11[47:0]  ), //i
    .Scale_dataIn_12  (bias_1_Bias_dataOut_12[47:0]  ), //i
    .Scale_dataIn_13  (bias_1_Bias_dataOut_13[47:0]  ), //i
    .Scale_dataIn_14  (bias_1_Bias_dataOut_14[47:0]  ), //i
    .Scale_dataIn_15  (bias_1_Bias_dataOut_15[47:0]  ), //i
    .Scale_quan_0     (_zz_Scale_quan_0_1[31:0]      ), //i
    .Scale_quan_1     (_zz_Scale_quan_1_1[31:0]      ), //i
    .Scale_quan_2     (_zz_Scale_quan_2_1[31:0]      ), //i
    .Scale_quan_3     (_zz_Scale_quan_3_1[31:0]      ), //i
    .Scale_quan_4     (_zz_Scale_quan_4_1[31:0]      ), //i
    .Scale_quan_5     (_zz_Scale_quan_5_1[31:0]      ), //i
    .Scale_quan_6     (_zz_Scale_quan_6_1[31:0]      ), //i
    .Scale_quan_7     (_zz_Scale_quan_7_1[31:0]      ), //i
    .Scale_quan_8     (_zz_Scale_quan_8_1[31:0]      ), //i
    .Scale_quan_9     (_zz_Scale_quan_9_1[31:0]      ), //i
    .Scale_quan_10    (_zz_Scale_quan_10_1[31:0]     ), //i
    .Scale_quan_11    (_zz_Scale_quan_11_1[31:0]     ), //i
    .Scale_quan_12    (_zz_Scale_quan_12_1[31:0]     ), //i
    .Scale_quan_13    (_zz_Scale_quan_13_1[31:0]     ), //i
    .Scale_quan_14    (_zz_Scale_quan_14_1[31:0]     ), //i
    .Scale_quan_15    (_zz_Scale_quan_15_1[31:0]     ), //i
    .Scale_dataOut_0  (scale_1_Scale_dataOut_0[31:0] ), //o
    .Scale_dataOut_1  (scale_1_Scale_dataOut_1[31:0] ), //o
    .Scale_dataOut_2  (scale_1_Scale_dataOut_2[31:0] ), //o
    .Scale_dataOut_3  (scale_1_Scale_dataOut_3[31:0] ), //o
    .Scale_dataOut_4  (scale_1_Scale_dataOut_4[31:0] ), //o
    .Scale_dataOut_5  (scale_1_Scale_dataOut_5[31:0] ), //o
    .Scale_dataOut_6  (scale_1_Scale_dataOut_6[31:0] ), //o
    .Scale_dataOut_7  (scale_1_Scale_dataOut_7[31:0] ), //o
    .Scale_dataOut_8  (scale_1_Scale_dataOut_8[31:0] ), //o
    .Scale_dataOut_9  (scale_1_Scale_dataOut_9[31:0] ), //o
    .Scale_dataOut_10 (scale_1_Scale_dataOut_10[31:0]), //o
    .Scale_dataOut_11 (scale_1_Scale_dataOut_11[31:0]), //o
    .Scale_dataOut_12 (scale_1_Scale_dataOut_12[31:0]), //o
    .Scale_dataOut_13 (scale_1_Scale_dataOut_13[31:0]), //o
    .Scale_dataOut_14 (scale_1_Scale_dataOut_14[31:0]), //o
    .Scale_dataOut_15 (scale_1_Scale_dataOut_15[31:0]), //o
    .clk              (clk                           ), //i
    .reset            (reset                         ), //i
    .softReset        (softReset                     )  //i
  );
  Shift shift_1 (
    .shift_dataIn_0   (scale_1_Scale_dataOut_0[31:0] ), //i
    .shift_dataIn_1   (scale_1_Scale_dataOut_1[31:0] ), //i
    .shift_dataIn_2   (scale_1_Scale_dataOut_2[31:0] ), //i
    .shift_dataIn_3   (scale_1_Scale_dataOut_3[31:0] ), //i
    .shift_dataIn_4   (scale_1_Scale_dataOut_4[31:0] ), //i
    .shift_dataIn_5   (scale_1_Scale_dataOut_5[31:0] ), //i
    .shift_dataIn_6   (scale_1_Scale_dataOut_6[31:0] ), //i
    .shift_dataIn_7   (scale_1_Scale_dataOut_7[31:0] ), //i
    .shift_dataIn_8   (scale_1_Scale_dataOut_8[31:0] ), //i
    .shift_dataIn_9   (scale_1_Scale_dataOut_9[31:0] ), //i
    .shift_dataIn_10  (scale_1_Scale_dataOut_10[31:0]), //i
    .shift_dataIn_11  (scale_1_Scale_dataOut_11[31:0]), //i
    .shift_dataIn_12  (scale_1_Scale_dataOut_12[31:0]), //i
    .shift_dataIn_13  (scale_1_Scale_dataOut_13[31:0]), //i
    .shift_dataIn_14  (scale_1_Scale_dataOut_14[31:0]), //i
    .shift_dataIn_15  (scale_1_Scale_dataOut_15[31:0]), //i
    .shift_quan_0     (_zz_shift_quan_0_10[31:0]     ), //i
    .shift_quan_1     (_zz_shift_quan_1_10[31:0]     ), //i
    .shift_quan_2     (_zz_shift_quan_2_10[31:0]     ), //i
    .shift_quan_3     (_zz_shift_quan_3_10[31:0]     ), //i
    .shift_quan_4     (_zz_shift_quan_4_10[31:0]     ), //i
    .shift_quan_5     (_zz_shift_quan_5_10[31:0]     ), //i
    .shift_quan_6     (_zz_shift_quan_6_10[31:0]     ), //i
    .shift_quan_7     (_zz_shift_quan_7_10[31:0]     ), //i
    .shift_quan_8     (_zz_shift_quan_8_10[31:0]     ), //i
    .shift_quan_9     (_zz_shift_quan_9_10[31:0]     ), //i
    .shift_quan_10    (_zz_shift_quan_10_10[31:0]    ), //i
    .shift_quan_11    (_zz_shift_quan_11_10[31:0]    ), //i
    .shift_quan_12    (_zz_shift_quan_12_10[31:0]    ), //i
    .shift_quan_13    (_zz_shift_quan_13_10[31:0]    ), //i
    .shift_quan_14    (_zz_shift_quan_14_10[31:0]    ), //i
    .shift_quan_15    (_zz_shift_quan_15_10[31:0]    ), //i
    .shift_dataOut_0  (shift_1_shift_dataOut_0[15:0] ), //o
    .shift_dataOut_1  (shift_1_shift_dataOut_1[15:0] ), //o
    .shift_dataOut_2  (shift_1_shift_dataOut_2[15:0] ), //o
    .shift_dataOut_3  (shift_1_shift_dataOut_3[15:0] ), //o
    .shift_dataOut_4  (shift_1_shift_dataOut_4[15:0] ), //o
    .shift_dataOut_5  (shift_1_shift_dataOut_5[15:0] ), //o
    .shift_dataOut_6  (shift_1_shift_dataOut_6[15:0] ), //o
    .shift_dataOut_7  (shift_1_shift_dataOut_7[15:0] ), //o
    .shift_dataOut_8  (shift_1_shift_dataOut_8[15:0] ), //o
    .shift_dataOut_9  (shift_1_shift_dataOut_9[15:0] ), //o
    .shift_dataOut_10 (shift_1_shift_dataOut_10[15:0]), //o
    .shift_dataOut_11 (shift_1_shift_dataOut_11[15:0]), //o
    .shift_dataOut_12 (shift_1_shift_dataOut_12[15:0]), //o
    .shift_dataOut_13 (shift_1_shift_dataOut_13[15:0]), //o
    .shift_dataOut_14 (shift_1_shift_dataOut_14[15:0]), //o
    .shift_dataOut_15 (shift_1_shift_dataOut_15[15:0]), //o
    .clk              (clk                           ), //i
    .reset            (reset                         ), //i
    .softReset        (softReset                     )  //i
  );
  Zero zero_1 (
    .dataIn_0   (shift_1_shift_dataOut_0[15:0] ), //i
    .dataIn_1   (shift_1_shift_dataOut_1[15:0] ), //i
    .dataIn_2   (shift_1_shift_dataOut_2[15:0] ), //i
    .dataIn_3   (shift_1_shift_dataOut_3[15:0] ), //i
    .dataIn_4   (shift_1_shift_dataOut_4[15:0] ), //i
    .dataIn_5   (shift_1_shift_dataOut_5[15:0] ), //i
    .dataIn_6   (shift_1_shift_dataOut_6[15:0] ), //i
    .dataIn_7   (shift_1_shift_dataOut_7[15:0] ), //i
    .dataIn_8   (shift_1_shift_dataOut_8[15:0] ), //i
    .dataIn_9   (shift_1_shift_dataOut_9[15:0] ), //i
    .dataIn_10  (shift_1_shift_dataOut_10[15:0]), //i
    .dataIn_11  (shift_1_shift_dataOut_11[15:0]), //i
    .dataIn_12  (shift_1_shift_dataOut_12[15:0]), //i
    .dataIn_13  (shift_1_shift_dataOut_13[15:0]), //i
    .dataIn_14  (shift_1_shift_dataOut_14[15:0]), //i
    .dataIn_15  (shift_1_shift_dataOut_15[15:0]), //i
    .quan_1     (zeroIn[7:0]                   ), //i
    .dataOut_0  (zero_1_dataOut_0[7:0]         ), //o
    .dataOut_1  (zero_1_dataOut_1[7:0]         ), //o
    .dataOut_2  (zero_1_dataOut_2[7:0]         ), //o
    .dataOut_3  (zero_1_dataOut_3[7:0]         ), //o
    .dataOut_4  (zero_1_dataOut_4[7:0]         ), //o
    .dataOut_5  (zero_1_dataOut_5[7:0]         ), //o
    .dataOut_6  (zero_1_dataOut_6[7:0]         ), //o
    .dataOut_7  (zero_1_dataOut_7[7:0]         ), //o
    .dataOut_8  (zero_1_dataOut_8[7:0]         ), //o
    .dataOut_9  (zero_1_dataOut_9[7:0]         ), //o
    .dataOut_10 (zero_1_dataOut_10[7:0]        ), //o
    .dataOut_11 (zero_1_dataOut_11[7:0]        ), //o
    .dataOut_12 (zero_1_dataOut_12[7:0]        ), //o
    .dataOut_13 (zero_1_dataOut_13[7:0]        ), //o
    .dataOut_14 (zero_1_dataOut_14[7:0]        ), //o
    .dataOut_15 (zero_1_dataOut_15[7:0]        ), //o
    .clk        (clk                           ), //i
    .reset      (reset                         ), //i
    .softReset  (softReset                     )  //i
  );
  LeakyRelu leakyRelu_1 (
    .dataIn_0   (zero_1_dataOut_0[7:0]      ), //i
    .dataIn_1   (zero_1_dataOut_1[7:0]      ), //i
    .dataIn_2   (zero_1_dataOut_2[7:0]      ), //i
    .dataIn_3   (zero_1_dataOut_3[7:0]      ), //i
    .dataIn_4   (zero_1_dataOut_4[7:0]      ), //i
    .dataIn_5   (zero_1_dataOut_5[7:0]      ), //i
    .dataIn_6   (zero_1_dataOut_6[7:0]      ), //i
    .dataIn_7   (zero_1_dataOut_7[7:0]      ), //i
    .dataIn_8   (zero_1_dataOut_8[7:0]      ), //i
    .dataIn_9   (zero_1_dataOut_9[7:0]      ), //i
    .dataIn_10  (zero_1_dataOut_10[7:0]     ), //i
    .dataIn_11  (zero_1_dataOut_11[7:0]     ), //i
    .dataIn_12  (zero_1_dataOut_12[7:0]     ), //i
    .dataIn_13  (zero_1_dataOut_13[7:0]     ), //i
    .dataIn_14  (zero_1_dataOut_14[7:0]     ), //i
    .dataIn_15  (zero_1_dataOut_15[7:0]     ), //i
    .quanZero   (zeroIn[7:0]                ), //i
    .amendReg   (amendReg[31:0]             ), //i
    .dataOut_0  (leakyRelu_1_dataOut_0[7:0] ), //o
    .dataOut_1  (leakyRelu_1_dataOut_1[7:0] ), //o
    .dataOut_2  (leakyRelu_1_dataOut_2[7:0] ), //o
    .dataOut_3  (leakyRelu_1_dataOut_3[7:0] ), //o
    .dataOut_4  (leakyRelu_1_dataOut_4[7:0] ), //o
    .dataOut_5  (leakyRelu_1_dataOut_5[7:0] ), //o
    .dataOut_6  (leakyRelu_1_dataOut_6[7:0] ), //o
    .dataOut_7  (leakyRelu_1_dataOut_7[7:0] ), //o
    .dataOut_8  (leakyRelu_1_dataOut_8[7:0] ), //o
    .dataOut_9  (leakyRelu_1_dataOut_9[7:0] ), //o
    .dataOut_10 (leakyRelu_1_dataOut_10[7:0]), //o
    .dataOut_11 (leakyRelu_1_dataOut_11[7:0]), //o
    .dataOut_12 (leakyRelu_1_dataOut_12[7:0]), //o
    .dataOut_13 (leakyRelu_1_dataOut_13[7:0]), //o
    .dataOut_14 (leakyRelu_1_dataOut_14[7:0]), //o
    .dataOut_15 (leakyRelu_1_dataOut_15[7:0]), //o
    .clk        (clk                        ), //i
    .reset      (reset                      ), //i
    .softReset  (softReset                  )  //i
  );
  assign bias_1_Bias_quan_0 = biasIn[31 : 0];
  assign bias_1_Bias_quan_1 = biasIn[63 : 32];
  assign bias_1_Bias_quan_2 = biasIn[95 : 64];
  assign bias_1_Bias_quan_3 = biasIn[127 : 96];
  assign bias_1_Bias_quan_4 = biasIn[159 : 128];
  assign bias_1_Bias_quan_5 = biasIn[191 : 160];
  assign bias_1_Bias_quan_6 = biasIn[223 : 192];
  assign bias_1_Bias_quan_7 = biasIn[255 : 224];
  assign bias_1_Bias_quan_8 = biasIn[287 : 256];
  assign bias_1_Bias_quan_9 = biasIn[319 : 288];
  assign bias_1_Bias_quan_10 = biasIn[351 : 320];
  assign bias_1_Bias_quan_11 = biasIn[383 : 352];
  assign bias_1_Bias_quan_12 = biasIn[415 : 384];
  assign bias_1_Bias_quan_13 = biasIn[447 : 416];
  assign bias_1_Bias_quan_14 = biasIn[479 : 448];
  assign bias_1_Bias_quan_15 = biasIn[511 : 480];
  always @(*) begin
    if(activationEn) begin
      dataOut[7 : 0] = leakyRelu_1_dataOut_0;
      dataOut[15 : 8] = leakyRelu_1_dataOut_1;
      dataOut[23 : 16] = leakyRelu_1_dataOut_2;
      dataOut[31 : 24] = leakyRelu_1_dataOut_3;
      dataOut[39 : 32] = leakyRelu_1_dataOut_4;
      dataOut[47 : 40] = leakyRelu_1_dataOut_5;
      dataOut[55 : 48] = leakyRelu_1_dataOut_6;
      dataOut[63 : 56] = leakyRelu_1_dataOut_7;
      dataOut[71 : 64] = leakyRelu_1_dataOut_8;
      dataOut[79 : 72] = leakyRelu_1_dataOut_9;
      dataOut[87 : 80] = leakyRelu_1_dataOut_10;
      dataOut[95 : 88] = leakyRelu_1_dataOut_11;
      dataOut[103 : 96] = leakyRelu_1_dataOut_12;
      dataOut[111 : 104] = leakyRelu_1_dataOut_13;
      dataOut[119 : 112] = leakyRelu_1_dataOut_14;
      dataOut[127 : 120] = leakyRelu_1_dataOut_15;
    end else begin
      dataOut[7 : 0] = zero_1_dataOut_0;
      dataOut[15 : 8] = zero_1_dataOut_1;
      dataOut[23 : 16] = zero_1_dataOut_2;
      dataOut[31 : 24] = zero_1_dataOut_3;
      dataOut[39 : 32] = zero_1_dataOut_4;
      dataOut[47 : 40] = zero_1_dataOut_5;
      dataOut[55 : 48] = zero_1_dataOut_6;
      dataOut[63 : 56] = zero_1_dataOut_7;
      dataOut[71 : 64] = zero_1_dataOut_8;
      dataOut[79 : 72] = zero_1_dataOut_9;
      dataOut[87 : 80] = zero_1_dataOut_10;
      dataOut[95 : 88] = zero_1_dataOut_11;
      dataOut[103 : 96] = zero_1_dataOut_12;
      dataOut[111 : 104] = zero_1_dataOut_13;
      dataOut[119 : 112] = zero_1_dataOut_14;
      dataOut[127 : 120] = zero_1_dataOut_15;
    end
  end

  always @(posedge clk) begin
    dataIn_regNext_0 <= dataIn_0;
    dataIn_regNext_1 <= dataIn_1;
    dataIn_regNext_2 <= dataIn_2;
    dataIn_regNext_3 <= dataIn_3;
    dataIn_regNext_4 <= dataIn_4;
    dataIn_regNext_5 <= dataIn_5;
    dataIn_regNext_6 <= dataIn_6;
    dataIn_regNext_7 <= dataIn_7;
    dataIn_regNext_8 <= dataIn_8;
    dataIn_regNext_9 <= dataIn_9;
    dataIn_regNext_10 <= dataIn_10;
    dataIn_regNext_11 <= dataIn_11;
    dataIn_regNext_12 <= dataIn_12;
    dataIn_regNext_13 <= dataIn_13;
    dataIn_regNext_14 <= dataIn_14;
    dataIn_regNext_15 <= dataIn_15;
    _zz_Scale_quan_0 <= scaleIn[31 : 0];
    _zz_Scale_quan_1 <= scaleIn[63 : 32];
    _zz_Scale_quan_2 <= scaleIn[95 : 64];
    _zz_Scale_quan_3 <= scaleIn[127 : 96];
    _zz_Scale_quan_4 <= scaleIn[159 : 128];
    _zz_Scale_quan_5 <= scaleIn[191 : 160];
    _zz_Scale_quan_6 <= scaleIn[223 : 192];
    _zz_Scale_quan_7 <= scaleIn[255 : 224];
    _zz_Scale_quan_8 <= scaleIn[287 : 256];
    _zz_Scale_quan_9 <= scaleIn[319 : 288];
    _zz_Scale_quan_10 <= scaleIn[351 : 320];
    _zz_Scale_quan_11 <= scaleIn[383 : 352];
    _zz_Scale_quan_12 <= scaleIn[415 : 384];
    _zz_Scale_quan_13 <= scaleIn[447 : 416];
    _zz_Scale_quan_14 <= scaleIn[479 : 448];
    _zz_Scale_quan_15 <= scaleIn[511 : 480];
    _zz_Scale_quan_0_1 <= _zz_Scale_quan_0;
    _zz_Scale_quan_1_1 <= _zz_Scale_quan_1;
    _zz_Scale_quan_2_1 <= _zz_Scale_quan_2;
    _zz_Scale_quan_3_1 <= _zz_Scale_quan_3;
    _zz_Scale_quan_4_1 <= _zz_Scale_quan_4;
    _zz_Scale_quan_5_1 <= _zz_Scale_quan_5;
    _zz_Scale_quan_6_1 <= _zz_Scale_quan_6;
    _zz_Scale_quan_7_1 <= _zz_Scale_quan_7;
    _zz_Scale_quan_8_1 <= _zz_Scale_quan_8;
    _zz_Scale_quan_9_1 <= _zz_Scale_quan_9;
    _zz_Scale_quan_10_1 <= _zz_Scale_quan_10;
    _zz_Scale_quan_11_1 <= _zz_Scale_quan_11;
    _zz_Scale_quan_12_1 <= _zz_Scale_quan_12;
    _zz_Scale_quan_13_1 <= _zz_Scale_quan_13;
    _zz_Scale_quan_14_1 <= _zz_Scale_quan_14;
    _zz_Scale_quan_15_1 <= _zz_Scale_quan_15;
    _zz_shift_quan_0 <= shiftIn[31 : 0];
    _zz_shift_quan_1 <= shiftIn[63 : 32];
    _zz_shift_quan_2 <= shiftIn[95 : 64];
    _zz_shift_quan_3 <= shiftIn[127 : 96];
    _zz_shift_quan_4 <= shiftIn[159 : 128];
    _zz_shift_quan_5 <= shiftIn[191 : 160];
    _zz_shift_quan_6 <= shiftIn[223 : 192];
    _zz_shift_quan_7 <= shiftIn[255 : 224];
    _zz_shift_quan_8 <= shiftIn[287 : 256];
    _zz_shift_quan_9 <= shiftIn[319 : 288];
    _zz_shift_quan_10 <= shiftIn[351 : 320];
    _zz_shift_quan_11 <= shiftIn[383 : 352];
    _zz_shift_quan_12 <= shiftIn[415 : 384];
    _zz_shift_quan_13 <= shiftIn[447 : 416];
    _zz_shift_quan_14 <= shiftIn[479 : 448];
    _zz_shift_quan_15 <= shiftIn[511 : 480];
    _zz_shift_quan_0_1 <= _zz_shift_quan_0;
    _zz_shift_quan_1_1 <= _zz_shift_quan_1;
    _zz_shift_quan_2_1 <= _zz_shift_quan_2;
    _zz_shift_quan_3_1 <= _zz_shift_quan_3;
    _zz_shift_quan_4_1 <= _zz_shift_quan_4;
    _zz_shift_quan_5_1 <= _zz_shift_quan_5;
    _zz_shift_quan_6_1 <= _zz_shift_quan_6;
    _zz_shift_quan_7_1 <= _zz_shift_quan_7;
    _zz_shift_quan_8_1 <= _zz_shift_quan_8;
    _zz_shift_quan_9_1 <= _zz_shift_quan_9;
    _zz_shift_quan_10_1 <= _zz_shift_quan_10;
    _zz_shift_quan_11_1 <= _zz_shift_quan_11;
    _zz_shift_quan_12_1 <= _zz_shift_quan_12;
    _zz_shift_quan_13_1 <= _zz_shift_quan_13;
    _zz_shift_quan_14_1 <= _zz_shift_quan_14;
    _zz_shift_quan_15_1 <= _zz_shift_quan_15;
    _zz_shift_quan_0_2 <= _zz_shift_quan_0_1;
    _zz_shift_quan_1_2 <= _zz_shift_quan_1_1;
    _zz_shift_quan_2_2 <= _zz_shift_quan_2_1;
    _zz_shift_quan_3_2 <= _zz_shift_quan_3_1;
    _zz_shift_quan_4_2 <= _zz_shift_quan_4_1;
    _zz_shift_quan_5_2 <= _zz_shift_quan_5_1;
    _zz_shift_quan_6_2 <= _zz_shift_quan_6_1;
    _zz_shift_quan_7_2 <= _zz_shift_quan_7_1;
    _zz_shift_quan_8_2 <= _zz_shift_quan_8_1;
    _zz_shift_quan_9_2 <= _zz_shift_quan_9_1;
    _zz_shift_quan_10_2 <= _zz_shift_quan_10_1;
    _zz_shift_quan_11_2 <= _zz_shift_quan_11_1;
    _zz_shift_quan_12_2 <= _zz_shift_quan_12_1;
    _zz_shift_quan_13_2 <= _zz_shift_quan_13_1;
    _zz_shift_quan_14_2 <= _zz_shift_quan_14_1;
    _zz_shift_quan_15_2 <= _zz_shift_quan_15_1;
    _zz_shift_quan_0_3 <= _zz_shift_quan_0_2;
    _zz_shift_quan_1_3 <= _zz_shift_quan_1_2;
    _zz_shift_quan_2_3 <= _zz_shift_quan_2_2;
    _zz_shift_quan_3_3 <= _zz_shift_quan_3_2;
    _zz_shift_quan_4_3 <= _zz_shift_quan_4_2;
    _zz_shift_quan_5_3 <= _zz_shift_quan_5_2;
    _zz_shift_quan_6_3 <= _zz_shift_quan_6_2;
    _zz_shift_quan_7_3 <= _zz_shift_quan_7_2;
    _zz_shift_quan_8_3 <= _zz_shift_quan_8_2;
    _zz_shift_quan_9_3 <= _zz_shift_quan_9_2;
    _zz_shift_quan_10_3 <= _zz_shift_quan_10_2;
    _zz_shift_quan_11_3 <= _zz_shift_quan_11_2;
    _zz_shift_quan_12_3 <= _zz_shift_quan_12_2;
    _zz_shift_quan_13_3 <= _zz_shift_quan_13_2;
    _zz_shift_quan_14_3 <= _zz_shift_quan_14_2;
    _zz_shift_quan_15_3 <= _zz_shift_quan_15_2;
    _zz_shift_quan_0_4 <= _zz_shift_quan_0_3;
    _zz_shift_quan_1_4 <= _zz_shift_quan_1_3;
    _zz_shift_quan_2_4 <= _zz_shift_quan_2_3;
    _zz_shift_quan_3_4 <= _zz_shift_quan_3_3;
    _zz_shift_quan_4_4 <= _zz_shift_quan_4_3;
    _zz_shift_quan_5_4 <= _zz_shift_quan_5_3;
    _zz_shift_quan_6_4 <= _zz_shift_quan_6_3;
    _zz_shift_quan_7_4 <= _zz_shift_quan_7_3;
    _zz_shift_quan_8_4 <= _zz_shift_quan_8_3;
    _zz_shift_quan_9_4 <= _zz_shift_quan_9_3;
    _zz_shift_quan_10_4 <= _zz_shift_quan_10_3;
    _zz_shift_quan_11_4 <= _zz_shift_quan_11_3;
    _zz_shift_quan_12_4 <= _zz_shift_quan_12_3;
    _zz_shift_quan_13_4 <= _zz_shift_quan_13_3;
    _zz_shift_quan_14_4 <= _zz_shift_quan_14_3;
    _zz_shift_quan_15_4 <= _zz_shift_quan_15_3;
    _zz_shift_quan_0_5 <= _zz_shift_quan_0_4;
    _zz_shift_quan_1_5 <= _zz_shift_quan_1_4;
    _zz_shift_quan_2_5 <= _zz_shift_quan_2_4;
    _zz_shift_quan_3_5 <= _zz_shift_quan_3_4;
    _zz_shift_quan_4_5 <= _zz_shift_quan_4_4;
    _zz_shift_quan_5_5 <= _zz_shift_quan_5_4;
    _zz_shift_quan_6_5 <= _zz_shift_quan_6_4;
    _zz_shift_quan_7_5 <= _zz_shift_quan_7_4;
    _zz_shift_quan_8_5 <= _zz_shift_quan_8_4;
    _zz_shift_quan_9_5 <= _zz_shift_quan_9_4;
    _zz_shift_quan_10_5 <= _zz_shift_quan_10_4;
    _zz_shift_quan_11_5 <= _zz_shift_quan_11_4;
    _zz_shift_quan_12_5 <= _zz_shift_quan_12_4;
    _zz_shift_quan_13_5 <= _zz_shift_quan_13_4;
    _zz_shift_quan_14_5 <= _zz_shift_quan_14_4;
    _zz_shift_quan_15_5 <= _zz_shift_quan_15_4;
    _zz_shift_quan_0_6 <= _zz_shift_quan_0_5;
    _zz_shift_quan_1_6 <= _zz_shift_quan_1_5;
    _zz_shift_quan_2_6 <= _zz_shift_quan_2_5;
    _zz_shift_quan_3_6 <= _zz_shift_quan_3_5;
    _zz_shift_quan_4_6 <= _zz_shift_quan_4_5;
    _zz_shift_quan_5_6 <= _zz_shift_quan_5_5;
    _zz_shift_quan_6_6 <= _zz_shift_quan_6_5;
    _zz_shift_quan_7_6 <= _zz_shift_quan_7_5;
    _zz_shift_quan_8_6 <= _zz_shift_quan_8_5;
    _zz_shift_quan_9_6 <= _zz_shift_quan_9_5;
    _zz_shift_quan_10_6 <= _zz_shift_quan_10_5;
    _zz_shift_quan_11_6 <= _zz_shift_quan_11_5;
    _zz_shift_quan_12_6 <= _zz_shift_quan_12_5;
    _zz_shift_quan_13_6 <= _zz_shift_quan_13_5;
    _zz_shift_quan_14_6 <= _zz_shift_quan_14_5;
    _zz_shift_quan_15_6 <= _zz_shift_quan_15_5;
    _zz_shift_quan_0_7 <= _zz_shift_quan_0_6;
    _zz_shift_quan_1_7 <= _zz_shift_quan_1_6;
    _zz_shift_quan_2_7 <= _zz_shift_quan_2_6;
    _zz_shift_quan_3_7 <= _zz_shift_quan_3_6;
    _zz_shift_quan_4_7 <= _zz_shift_quan_4_6;
    _zz_shift_quan_5_7 <= _zz_shift_quan_5_6;
    _zz_shift_quan_6_7 <= _zz_shift_quan_6_6;
    _zz_shift_quan_7_7 <= _zz_shift_quan_7_6;
    _zz_shift_quan_8_7 <= _zz_shift_quan_8_6;
    _zz_shift_quan_9_7 <= _zz_shift_quan_9_6;
    _zz_shift_quan_10_7 <= _zz_shift_quan_10_6;
    _zz_shift_quan_11_7 <= _zz_shift_quan_11_6;
    _zz_shift_quan_12_7 <= _zz_shift_quan_12_6;
    _zz_shift_quan_13_7 <= _zz_shift_quan_13_6;
    _zz_shift_quan_14_7 <= _zz_shift_quan_14_6;
    _zz_shift_quan_15_7 <= _zz_shift_quan_15_6;
    _zz_shift_quan_0_8 <= _zz_shift_quan_0_7;
    _zz_shift_quan_1_8 <= _zz_shift_quan_1_7;
    _zz_shift_quan_2_8 <= _zz_shift_quan_2_7;
    _zz_shift_quan_3_8 <= _zz_shift_quan_3_7;
    _zz_shift_quan_4_8 <= _zz_shift_quan_4_7;
    _zz_shift_quan_5_8 <= _zz_shift_quan_5_7;
    _zz_shift_quan_6_8 <= _zz_shift_quan_6_7;
    _zz_shift_quan_7_8 <= _zz_shift_quan_7_7;
    _zz_shift_quan_8_8 <= _zz_shift_quan_8_7;
    _zz_shift_quan_9_8 <= _zz_shift_quan_9_7;
    _zz_shift_quan_10_8 <= _zz_shift_quan_10_7;
    _zz_shift_quan_11_8 <= _zz_shift_quan_11_7;
    _zz_shift_quan_12_8 <= _zz_shift_quan_12_7;
    _zz_shift_quan_13_8 <= _zz_shift_quan_13_7;
    _zz_shift_quan_14_8 <= _zz_shift_quan_14_7;
    _zz_shift_quan_15_8 <= _zz_shift_quan_15_7;
    _zz_shift_quan_0_9 <= _zz_shift_quan_0_8;
    _zz_shift_quan_1_9 <= _zz_shift_quan_1_8;
    _zz_shift_quan_2_9 <= _zz_shift_quan_2_8;
    _zz_shift_quan_3_9 <= _zz_shift_quan_3_8;
    _zz_shift_quan_4_9 <= _zz_shift_quan_4_8;
    _zz_shift_quan_5_9 <= _zz_shift_quan_5_8;
    _zz_shift_quan_6_9 <= _zz_shift_quan_6_8;
    _zz_shift_quan_7_9 <= _zz_shift_quan_7_8;
    _zz_shift_quan_8_9 <= _zz_shift_quan_8_8;
    _zz_shift_quan_9_9 <= _zz_shift_quan_9_8;
    _zz_shift_quan_10_9 <= _zz_shift_quan_10_8;
    _zz_shift_quan_11_9 <= _zz_shift_quan_11_8;
    _zz_shift_quan_12_9 <= _zz_shift_quan_12_8;
    _zz_shift_quan_13_9 <= _zz_shift_quan_13_8;
    _zz_shift_quan_14_9 <= _zz_shift_quan_14_8;
    _zz_shift_quan_15_9 <= _zz_shift_quan_15_8;
    _zz_shift_quan_0_10 <= _zz_shift_quan_0_9;
    _zz_shift_quan_1_10 <= _zz_shift_quan_1_9;
    _zz_shift_quan_2_10 <= _zz_shift_quan_2_9;
    _zz_shift_quan_3_10 <= _zz_shift_quan_3_9;
    _zz_shift_quan_4_10 <= _zz_shift_quan_4_9;
    _zz_shift_quan_5_10 <= _zz_shift_quan_5_9;
    _zz_shift_quan_6_10 <= _zz_shift_quan_6_9;
    _zz_shift_quan_7_10 <= _zz_shift_quan_7_9;
    _zz_shift_quan_8_10 <= _zz_shift_quan_8_9;
    _zz_shift_quan_9_10 <= _zz_shift_quan_9_9;
    _zz_shift_quan_10_10 <= _zz_shift_quan_10_9;
    _zz_shift_quan_11_10 <= _zz_shift_quan_11_9;
    _zz_shift_quan_12_10 <= _zz_shift_quan_12_9;
    _zz_shift_quan_13_10 <= _zz_shift_quan_13_9;
    _zz_shift_quan_14_10 <= _zz_shift_quan_14_9;
    _zz_shift_quan_15_10 <= _zz_shift_quan_15_9;
  end


endmodule

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

//xAddChannelTimes replaced by xAddChannelTimes

module xAddChannelTimes (
  input      [23:0]   A,
  output     [31:0]   S,
  input               init,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [31:0]   _zz_temp;
  reg        [31:0]   S_1;
  (* use_dsp = "yes" *) reg        [31:0]   temp;

  assign _zz_temp = {{8{A[23]}}, A};
  always @(*) begin
    if(init) begin
      S_1 = 32'h0;
    end else begin
      S_1 = temp;
    end
  end

  assign S = temp;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      temp <= 32'h0;
    end else begin
      if(softReset) begin
      temp <= 32'h0;
      end else begin
        temp <= ($signed(_zz_temp) + $signed(S_1));
      end
    end
  end


endmodule

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

//xAddTimes_128 replaced by xAddTimes_128

module xAddTimes_128 (
  input      [39:0]   A_0,
  input      [39:0]   A_1,
  input      [39:0]   A_2,
  input      [39:0]   A_3,
  input      [39:0]   A_4,
  input      [39:0]   A_5,
  input      [39:0]   A_6,
  input      [39:0]   A_7,
  input      [39:0]   A_8,
  input      [39:0]   A_9,
  input      [39:0]   A_10,
  input      [39:0]   A_11,
  input      [39:0]   A_12,
  input      [39:0]   A_13,
  input      [39:0]   A_14,
  input      [39:0]   A_15,
  output     [47:0]   S,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [20:0]   _zz__zz_S;
  wire       [20:0]   _zz__zz_S_1;
  wire       [20:0]   _zz__zz_S_1_1;
  wire       [20:0]   _zz__zz_S_1_2;
  wire       [20:0]   _zz__zz_S_2;
  wire       [20:0]   _zz__zz_S_2_1;
  wire       [20:0]   _zz__zz_S_3;
  wire       [20:0]   _zz__zz_S_3_1;
  wire       [20:0]   _zz__zz_S_4;
  wire       [20:0]   _zz__zz_S_4_1;
  wire       [20:0]   _zz__zz_S_5;
  wire       [20:0]   _zz__zz_S_5_1;
  wire       [20:0]   _zz__zz_S_6;
  wire       [20:0]   _zz__zz_S_6_1;
  wire       [20:0]   _zz__zz_S_7;
  wire       [20:0]   _zz__zz_S_7_1;
  wire       [21:0]   _zz__zz_S_8;
  wire       [21:0]   _zz__zz_S_8_1;
  wire       [21:0]   _zz__zz_S_9;
  wire       [21:0]   _zz__zz_S_9_1;
  wire       [21:0]   _zz__zz_S_10;
  wire       [21:0]   _zz__zz_S_10_1;
  wire       [21:0]   _zz__zz_S_11;
  wire       [21:0]   _zz__zz_S_11_1;
  wire       [22:0]   _zz__zz_S_12;
  wire       [22:0]   _zz__zz_S_12_1;
  wire       [22:0]   _zz__zz_S_13;
  wire       [22:0]   _zz__zz_S_13_1;
  wire       [23:0]   _zz__zz_S_14;
  wire       [23:0]   _zz__zz_S_14_1;
  wire       [20:0]   _zz__zz_S_15;
  wire       [20:0]   _zz__zz_S_15_1;
  wire       [20:0]   _zz__zz_S_16;
  wire       [20:0]   _zz__zz_S_16_1;
  wire       [20:0]   _zz__zz_S_17;
  wire       [20:0]   _zz__zz_S_17_1;
  wire       [20:0]   _zz__zz_S_18;
  wire       [20:0]   _zz__zz_S_18_1;
  wire       [20:0]   _zz__zz_S_19;
  wire       [20:0]   _zz__zz_S_19_1;
  wire       [20:0]   _zz__zz_S_20;
  wire       [20:0]   _zz__zz_S_20_1;
  wire       [20:0]   _zz__zz_S_21;
  wire       [20:0]   _zz__zz_S_21_1;
  wire       [20:0]   _zz__zz_S_22;
  wire       [20:0]   _zz__zz_S_22_1;
  wire       [21:0]   _zz__zz_S_23;
  wire       [21:0]   _zz__zz_S_23_1;
  wire       [21:0]   _zz__zz_S_24;
  wire       [21:0]   _zz__zz_S_24_1;
  wire       [21:0]   _zz__zz_S_25;
  wire       [21:0]   _zz__zz_S_25_1;
  wire       [21:0]   _zz__zz_S_26;
  wire       [21:0]   _zz__zz_S_26_1;
  wire       [22:0]   _zz__zz_S_27;
  wire       [22:0]   _zz__zz_S_27_1;
  wire       [22:0]   _zz__zz_S_28;
  wire       [22:0]   _zz__zz_S_28_1;
  wire       [23:0]   _zz__zz_S_29;
  wire       [23:0]   _zz__zz_S_29_1;
  wire       [19:0]   a1Temp_0;
  wire       [19:0]   a1Temp_1;
  wire       [19:0]   a1Temp_2;
  wire       [19:0]   a1Temp_3;
  wire       [19:0]   a1Temp_4;
  wire       [19:0]   a1Temp_5;
  wire       [19:0]   a1Temp_6;
  wire       [19:0]   a1Temp_7;
  wire       [19:0]   a1Temp_8;
  wire       [19:0]   a1Temp_9;
  wire       [19:0]   a1Temp_10;
  wire       [19:0]   a1Temp_11;
  wire       [19:0]   a1Temp_12;
  wire       [19:0]   a1Temp_13;
  wire       [19:0]   a1Temp_14;
  wire       [19:0]   a1Temp_15;
  wire       [19:0]   a2Temp_0;
  wire       [19:0]   a2Temp_1;
  wire       [19:0]   a2Temp_2;
  wire       [19:0]   a2Temp_3;
  wire       [19:0]   a2Temp_4;
  wire       [19:0]   a2Temp_5;
  wire       [19:0]   a2Temp_6;
  wire       [19:0]   a2Temp_7;
  wire       [19:0]   a2Temp_8;
  wire       [19:0]   a2Temp_9;
  wire       [19:0]   a2Temp_10;
  wire       [19:0]   a2Temp_11;
  wire       [19:0]   a2Temp_12;
  wire       [19:0]   a2Temp_13;
  wire       [19:0]   a2Temp_14;
  wire       [19:0]   a2Temp_15;
  reg        [20:0]   _zz_S;
  reg        [20:0]   _zz_S_1;
  reg        [20:0]   _zz_S_2;
  reg        [20:0]   _zz_S_3;
  reg        [20:0]   _zz_S_4;
  reg        [20:0]   _zz_S_5;
  reg        [20:0]   _zz_S_6;
  reg        [20:0]   _zz_S_7;
  reg        [21:0]   _zz_S_8;
  reg        [21:0]   _zz_S_9;
  reg        [21:0]   _zz_S_10;
  reg        [21:0]   _zz_S_11;
  reg        [22:0]   _zz_S_12;
  reg        [22:0]   _zz_S_13;
  reg        [23:0]   _zz_S_14;
  reg        [20:0]   _zz_S_15;
  reg        [20:0]   _zz_S_16;
  reg        [20:0]   _zz_S_17;
  reg        [20:0]   _zz_S_18;
  reg        [20:0]   _zz_S_19;
  reg        [20:0]   _zz_S_20;
  reg        [20:0]   _zz_S_21;
  reg        [20:0]   _zz_S_22;
  reg        [21:0]   _zz_S_23;
  reg        [21:0]   _zz_S_24;
  reg        [21:0]   _zz_S_25;
  reg        [21:0]   _zz_S_26;
  reg        [22:0]   _zz_S_27;
  reg        [22:0]   _zz_S_28;
  reg        [23:0]   _zz_S_29;

  assign _zz__zz_S = {a2Temp_0[19],a2Temp_0};
  assign _zz__zz_S_1 = {a2Temp_1[19],a2Temp_1};
  assign _zz__zz_S_1_1 = {a2Temp_2[19],a2Temp_2};
  assign _zz__zz_S_1_2 = {a2Temp_3[19],a2Temp_3};
  assign _zz__zz_S_2 = {a2Temp_4[19],a2Temp_4};
  assign _zz__zz_S_2_1 = {a2Temp_5[19],a2Temp_5};
  assign _zz__zz_S_3 = {a2Temp_6[19],a2Temp_6};
  assign _zz__zz_S_3_1 = {a2Temp_7[19],a2Temp_7};
  assign _zz__zz_S_4 = {a2Temp_8[19],a2Temp_8};
  assign _zz__zz_S_4_1 = {a2Temp_9[19],a2Temp_9};
  assign _zz__zz_S_5 = {a2Temp_10[19],a2Temp_10};
  assign _zz__zz_S_5_1 = {a2Temp_11[19],a2Temp_11};
  assign _zz__zz_S_6 = {a2Temp_12[19],a2Temp_12};
  assign _zz__zz_S_6_1 = {a2Temp_13[19],a2Temp_13};
  assign _zz__zz_S_7 = {a2Temp_14[19],a2Temp_14};
  assign _zz__zz_S_7_1 = {a2Temp_15[19],a2Temp_15};
  assign _zz__zz_S_8 = {_zz_S[20],_zz_S};
  assign _zz__zz_S_8_1 = {_zz_S_1[20],_zz_S_1};
  assign _zz__zz_S_9 = {_zz_S_2[20],_zz_S_2};
  assign _zz__zz_S_9_1 = {_zz_S_3[20],_zz_S_3};
  assign _zz__zz_S_10 = {_zz_S_4[20],_zz_S_4};
  assign _zz__zz_S_10_1 = {_zz_S_5[20],_zz_S_5};
  assign _zz__zz_S_11 = {_zz_S_6[20],_zz_S_6};
  assign _zz__zz_S_11_1 = {_zz_S_7[20],_zz_S_7};
  assign _zz__zz_S_12 = {_zz_S_8[21],_zz_S_8};
  assign _zz__zz_S_12_1 = {_zz_S_9[21],_zz_S_9};
  assign _zz__zz_S_13 = {_zz_S_10[21],_zz_S_10};
  assign _zz__zz_S_13_1 = {_zz_S_11[21],_zz_S_11};
  assign _zz__zz_S_14 = {_zz_S_12[22],_zz_S_12};
  assign _zz__zz_S_14_1 = {_zz_S_13[22],_zz_S_13};
  assign _zz__zz_S_15 = {a1Temp_0[19],a1Temp_0};
  assign _zz__zz_S_15_1 = {a1Temp_1[19],a1Temp_1};
  assign _zz__zz_S_16 = {a1Temp_2[19],a1Temp_2};
  assign _zz__zz_S_16_1 = {a1Temp_3[19],a1Temp_3};
  assign _zz__zz_S_17 = {a1Temp_4[19],a1Temp_4};
  assign _zz__zz_S_17_1 = {a1Temp_5[19],a1Temp_5};
  assign _zz__zz_S_18 = {a1Temp_6[19],a1Temp_6};
  assign _zz__zz_S_18_1 = {a1Temp_7[19],a1Temp_7};
  assign _zz__zz_S_19 = {a1Temp_8[19],a1Temp_8};
  assign _zz__zz_S_19_1 = {a1Temp_9[19],a1Temp_9};
  assign _zz__zz_S_20 = {a1Temp_10[19],a1Temp_10};
  assign _zz__zz_S_20_1 = {a1Temp_11[19],a1Temp_11};
  assign _zz__zz_S_21 = {a1Temp_12[19],a1Temp_12};
  assign _zz__zz_S_21_1 = {a1Temp_13[19],a1Temp_13};
  assign _zz__zz_S_22 = {a1Temp_14[19],a1Temp_14};
  assign _zz__zz_S_22_1 = {a1Temp_15[19],a1Temp_15};
  assign _zz__zz_S_23 = {_zz_S_15[20],_zz_S_15};
  assign _zz__zz_S_23_1 = {_zz_S_16[20],_zz_S_16};
  assign _zz__zz_S_24 = {_zz_S_17[20],_zz_S_17};
  assign _zz__zz_S_24_1 = {_zz_S_18[20],_zz_S_18};
  assign _zz__zz_S_25 = {_zz_S_19[20],_zz_S_19};
  assign _zz__zz_S_25_1 = {_zz_S_20[20],_zz_S_20};
  assign _zz__zz_S_26 = {_zz_S_21[20],_zz_S_21};
  assign _zz__zz_S_26_1 = {_zz_S_22[20],_zz_S_22};
  assign _zz__zz_S_27 = {_zz_S_23[21],_zz_S_23};
  assign _zz__zz_S_27_1 = {_zz_S_24[21],_zz_S_24};
  assign _zz__zz_S_28 = {_zz_S_25[21],_zz_S_25};
  assign _zz__zz_S_28_1 = {_zz_S_26[21],_zz_S_26};
  assign _zz__zz_S_29 = {_zz_S_27[22],_zz_S_27};
  assign _zz__zz_S_29_1 = {_zz_S_28[22],_zz_S_28};
  assign a1Temp_0 = A_0[19 : 0];
  assign a2Temp_0 = A_0[39 : 20];
  assign a1Temp_1 = A_1[19 : 0];
  assign a2Temp_1 = A_1[39 : 20];
  assign a1Temp_2 = A_2[19 : 0];
  assign a2Temp_2 = A_2[39 : 20];
  assign a1Temp_3 = A_3[19 : 0];
  assign a2Temp_3 = A_3[39 : 20];
  assign a1Temp_4 = A_4[19 : 0];
  assign a2Temp_4 = A_4[39 : 20];
  assign a1Temp_5 = A_5[19 : 0];
  assign a2Temp_5 = A_5[39 : 20];
  assign a1Temp_6 = A_6[19 : 0];
  assign a2Temp_6 = A_6[39 : 20];
  assign a1Temp_7 = A_7[19 : 0];
  assign a2Temp_7 = A_7[39 : 20];
  assign a1Temp_8 = A_8[19 : 0];
  assign a2Temp_8 = A_8[39 : 20];
  assign a1Temp_9 = A_9[19 : 0];
  assign a2Temp_9 = A_9[39 : 20];
  assign a1Temp_10 = A_10[19 : 0];
  assign a2Temp_10 = A_10[39 : 20];
  assign a1Temp_11 = A_11[19 : 0];
  assign a2Temp_11 = A_11[39 : 20];
  assign a1Temp_12 = A_12[19 : 0];
  assign a2Temp_12 = A_12[39 : 20];
  assign a1Temp_13 = A_13[19 : 0];
  assign a2Temp_13 = A_13[39 : 20];
  assign a1Temp_14 = A_14[19 : 0];
  assign a2Temp_14 = A_14[39 : 20];
  assign a1Temp_15 = A_15[19 : 0];
  assign a2Temp_15 = A_15[39 : 20];
  assign S = {_zz_S_14,_zz_S_29};
  always @(posedge clk) begin
    _zz_S <= ($signed(_zz__zz_S) + $signed(_zz__zz_S_1));
    _zz_S_1 <= ($signed(_zz__zz_S_1_1) + $signed(_zz__zz_S_1_2));
    _zz_S_2 <= ($signed(_zz__zz_S_2) + $signed(_zz__zz_S_2_1));
    _zz_S_3 <= ($signed(_zz__zz_S_3) + $signed(_zz__zz_S_3_1));
    _zz_S_4 <= ($signed(_zz__zz_S_4) + $signed(_zz__zz_S_4_1));
    _zz_S_5 <= ($signed(_zz__zz_S_5) + $signed(_zz__zz_S_5_1));
    _zz_S_6 <= ($signed(_zz__zz_S_6) + $signed(_zz__zz_S_6_1));
    _zz_S_7 <= ($signed(_zz__zz_S_7) + $signed(_zz__zz_S_7_1));
    _zz_S_8 <= ($signed(_zz__zz_S_8) + $signed(_zz__zz_S_8_1));
    _zz_S_9 <= ($signed(_zz__zz_S_9) + $signed(_zz__zz_S_9_1));
    _zz_S_10 <= ($signed(_zz__zz_S_10) + $signed(_zz__zz_S_10_1));
    _zz_S_11 <= ($signed(_zz__zz_S_11) + $signed(_zz__zz_S_11_1));
    _zz_S_12 <= ($signed(_zz__zz_S_12) + $signed(_zz__zz_S_12_1));
    _zz_S_13 <= ($signed(_zz__zz_S_13) + $signed(_zz__zz_S_13_1));
    _zz_S_14 <= ($signed(_zz__zz_S_14) + $signed(_zz__zz_S_14_1));
    _zz_S_15 <= ($signed(_zz__zz_S_15) + $signed(_zz__zz_S_15_1));
    _zz_S_16 <= ($signed(_zz__zz_S_16) + $signed(_zz__zz_S_16_1));
    _zz_S_17 <= ($signed(_zz__zz_S_17) + $signed(_zz__zz_S_17_1));
    _zz_S_18 <= ($signed(_zz__zz_S_18) + $signed(_zz__zz_S_18_1));
    _zz_S_19 <= ($signed(_zz__zz_S_19) + $signed(_zz__zz_S_19_1));
    _zz_S_20 <= ($signed(_zz__zz_S_20) + $signed(_zz__zz_S_20_1));
    _zz_S_21 <= ($signed(_zz__zz_S_21) + $signed(_zz__zz_S_21_1));
    _zz_S_22 <= ($signed(_zz__zz_S_22) + $signed(_zz__zz_S_22_1));
    _zz_S_23 <= ($signed(_zz__zz_S_23) + $signed(_zz__zz_S_23_1));
    _zz_S_24 <= ($signed(_zz__zz_S_24) + $signed(_zz__zz_S_24_1));
    _zz_S_25 <= ($signed(_zz__zz_S_25) + $signed(_zz__zz_S_25_1));
    _zz_S_26 <= ($signed(_zz__zz_S_26) + $signed(_zz__zz_S_26_1));
    _zz_S_27 <= ($signed(_zz__zz_S_27) + $signed(_zz__zz_S_27_1));
    _zz_S_28 <= ($signed(_zz__zz_S_28) + $signed(_zz__zz_S_28_1));
    _zz_S_29 <= ($signed(_zz__zz_S_29) + $signed(_zz__zz_S_29_1));
  end


endmodule

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

//xAddTimes replaced by xAddTimes

module xAddTimes (
  input      [31:0]   A_0,
  input      [31:0]   A_1,
  input      [31:0]   A_2,
  input      [31:0]   A_3,
  input      [31:0]   A_4,
  input      [31:0]   A_5,
  input      [31:0]   A_6,
  input      [31:0]   A_7,
  input      [31:0]   A_8,
  output     [39:0]   S,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [16:0]   _zz__zz_S;
  wire       [16:0]   _zz__zz_S_1;
  wire       [16:0]   _zz__zz_S_1_1;
  wire       [16:0]   _zz__zz_S_1_2;
  wire       [16:0]   _zz__zz_S_2;
  wire       [16:0]   _zz__zz_S_2_1;
  wire       [16:0]   _zz__zz_S_3;
  wire       [16:0]   _zz__zz_S_3_1;
  wire       [17:0]   _zz__zz_S_4;
  wire       [17:0]   _zz__zz_S_4_1;
  wire       [17:0]   _zz__zz_S_5;
  wire       [17:0]   _zz__zz_S_5_1;
  wire       [18:0]   _zz__zz_S_6;
  wire       [18:0]   _zz__zz_S_6_1;
  wire       [19:0]   _zz__zz_S_7;
  wire       [19:0]   _zz__zz_S_7_1;
  wire       [16:0]   _zz__zz_S_7_2;
  wire       [16:0]   _zz__zz_S_8;
  wire       [16:0]   _zz__zz_S_8_1;
  wire       [16:0]   _zz__zz_S_9;
  wire       [16:0]   _zz__zz_S_9_1;
  wire       [16:0]   _zz__zz_S_10;
  wire       [16:0]   _zz__zz_S_10_1;
  wire       [16:0]   _zz__zz_S_11;
  wire       [16:0]   _zz__zz_S_11_1;
  wire       [17:0]   _zz__zz_S_12;
  wire       [17:0]   _zz__zz_S_12_1;
  wire       [17:0]   _zz__zz_S_13;
  wire       [17:0]   _zz__zz_S_13_1;
  wire       [18:0]   _zz__zz_S_14;
  wire       [18:0]   _zz__zz_S_14_1;
  wire       [19:0]   _zz__zz_S_15;
  wire       [19:0]   _zz__zz_S_15_1;
  wire       [16:0]   _zz__zz_S_15_2;
  wire       [15:0]   a1Temp_0;
  wire       [15:0]   a1Temp_1;
  wire       [15:0]   a1Temp_2;
  wire       [15:0]   a1Temp_3;
  wire       [15:0]   a1Temp_4;
  wire       [15:0]   a1Temp_5;
  wire       [15:0]   a1Temp_6;
  wire       [15:0]   a1Temp_7;
  wire       [15:0]   a1Temp_8;
  wire       [15:0]   a2Temp_0;
  wire       [15:0]   a2Temp_1;
  wire       [15:0]   a2Temp_2;
  wire       [15:0]   a2Temp_3;
  wire       [15:0]   a2Temp_4;
  wire       [15:0]   a2Temp_5;
  wire       [15:0]   a2Temp_6;
  wire       [15:0]   a2Temp_7;
  wire       [15:0]   a2Temp_8;
  reg        [16:0]   _zz_S;
  reg        [16:0]   _zz_S_1;
  reg        [16:0]   _zz_S_2;
  reg        [16:0]   _zz_S_3;
  reg        [15:0]   a2Temp_8_regNext;
  reg        [17:0]   _zz_S_4;
  reg        [17:0]   _zz_S_5;
  reg        [15:0]   a2Temp_8_regNext_regNext;
  reg        [18:0]   _zz_S_6;
  reg        [15:0]   a2Temp_8_regNext_regNext_regNext;
  reg        [19:0]   _zz_S_7;
  reg        [16:0]   _zz_S_8;
  reg        [16:0]   _zz_S_9;
  reg        [16:0]   _zz_S_10;
  reg        [16:0]   _zz_S_11;
  reg        [15:0]   a1Temp_8_regNext;
  reg        [17:0]   _zz_S_12;
  reg        [17:0]   _zz_S_13;
  reg        [15:0]   a1Temp_8_regNext_regNext;
  reg        [18:0]   _zz_S_14;
  reg        [15:0]   a1Temp_8_regNext_regNext_regNext;
  reg        [19:0]   _zz_S_15;

  assign _zz__zz_S = {a2Temp_0[15],a2Temp_0};
  assign _zz__zz_S_1 = {a2Temp_1[15],a2Temp_1};
  assign _zz__zz_S_1_1 = {a2Temp_2[15],a2Temp_2};
  assign _zz__zz_S_1_2 = {a2Temp_3[15],a2Temp_3};
  assign _zz__zz_S_2 = {a2Temp_4[15],a2Temp_4};
  assign _zz__zz_S_2_1 = {a2Temp_5[15],a2Temp_5};
  assign _zz__zz_S_3 = {a2Temp_6[15],a2Temp_6};
  assign _zz__zz_S_3_1 = {a2Temp_7[15],a2Temp_7};
  assign _zz__zz_S_4 = {_zz_S[16],_zz_S};
  assign _zz__zz_S_4_1 = {_zz_S_1[16],_zz_S_1};
  assign _zz__zz_S_5 = {_zz_S_2[16],_zz_S_2};
  assign _zz__zz_S_5_1 = {_zz_S_3[16],_zz_S_3};
  assign _zz__zz_S_6 = {_zz_S_4[17],_zz_S_4};
  assign _zz__zz_S_6_1 = {_zz_S_5[17],_zz_S_5};
  assign _zz__zz_S_7 = {_zz_S_6[18],_zz_S_6};
  assign _zz__zz_S_7_2 = {a2Temp_8_regNext_regNext_regNext[15],a2Temp_8_regNext_regNext_regNext};
  assign _zz__zz_S_7_1 = {{3{_zz__zz_S_7_2[16]}}, _zz__zz_S_7_2};
  assign _zz__zz_S_8 = {a1Temp_0[15],a1Temp_0};
  assign _zz__zz_S_8_1 = {a1Temp_1[15],a1Temp_1};
  assign _zz__zz_S_9 = {a1Temp_2[15],a1Temp_2};
  assign _zz__zz_S_9_1 = {a1Temp_3[15],a1Temp_3};
  assign _zz__zz_S_10 = {a1Temp_4[15],a1Temp_4};
  assign _zz__zz_S_10_1 = {a1Temp_5[15],a1Temp_5};
  assign _zz__zz_S_11 = {a1Temp_6[15],a1Temp_6};
  assign _zz__zz_S_11_1 = {a1Temp_7[15],a1Temp_7};
  assign _zz__zz_S_12 = {_zz_S_8[16],_zz_S_8};
  assign _zz__zz_S_12_1 = {_zz_S_9[16],_zz_S_9};
  assign _zz__zz_S_13 = {_zz_S_10[16],_zz_S_10};
  assign _zz__zz_S_13_1 = {_zz_S_11[16],_zz_S_11};
  assign _zz__zz_S_14 = {_zz_S_12[17],_zz_S_12};
  assign _zz__zz_S_14_1 = {_zz_S_13[17],_zz_S_13};
  assign _zz__zz_S_15 = {_zz_S_14[18],_zz_S_14};
  assign _zz__zz_S_15_2 = {a1Temp_8_regNext_regNext_regNext[15],a1Temp_8_regNext_regNext_regNext};
  assign _zz__zz_S_15_1 = {{3{_zz__zz_S_15_2[16]}}, _zz__zz_S_15_2};
  assign a1Temp_0 = A_0[15 : 0];
  assign a2Temp_0 = A_0[31 : 16];
  assign a1Temp_1 = A_1[15 : 0];
  assign a2Temp_1 = A_1[31 : 16];
  assign a1Temp_2 = A_2[15 : 0];
  assign a2Temp_2 = A_2[31 : 16];
  assign a1Temp_3 = A_3[15 : 0];
  assign a2Temp_3 = A_3[31 : 16];
  assign a1Temp_4 = A_4[15 : 0];
  assign a2Temp_4 = A_4[31 : 16];
  assign a1Temp_5 = A_5[15 : 0];
  assign a2Temp_5 = A_5[31 : 16];
  assign a1Temp_6 = A_6[15 : 0];
  assign a2Temp_6 = A_6[31 : 16];
  assign a1Temp_7 = A_7[15 : 0];
  assign a2Temp_7 = A_7[31 : 16];
  assign a1Temp_8 = A_8[15 : 0];
  assign a2Temp_8 = A_8[31 : 16];
  assign S = {_zz_S_7,_zz_S_15};
  always @(posedge clk) begin
    _zz_S <= ($signed(_zz__zz_S) + $signed(_zz__zz_S_1));
    _zz_S_1 <= ($signed(_zz__zz_S_1_1) + $signed(_zz__zz_S_1_2));
    _zz_S_2 <= ($signed(_zz__zz_S_2) + $signed(_zz__zz_S_2_1));
    _zz_S_3 <= ($signed(_zz__zz_S_3) + $signed(_zz__zz_S_3_1));
    a2Temp_8_regNext <= a2Temp_8;
    _zz_S_4 <= ($signed(_zz__zz_S_4) + $signed(_zz__zz_S_4_1));
    _zz_S_5 <= ($signed(_zz__zz_S_5) + $signed(_zz__zz_S_5_1));
    a2Temp_8_regNext_regNext <= a2Temp_8_regNext;
    _zz_S_6 <= ($signed(_zz__zz_S_6) + $signed(_zz__zz_S_6_1));
    a2Temp_8_regNext_regNext_regNext <= a2Temp_8_regNext_regNext;
    _zz_S_7 <= ($signed(_zz__zz_S_7) + $signed(_zz__zz_S_7_1));
    _zz_S_8 <= ($signed(_zz__zz_S_8) + $signed(_zz__zz_S_8_1));
    _zz_S_9 <= ($signed(_zz__zz_S_9) + $signed(_zz__zz_S_9_1));
    _zz_S_10 <= ($signed(_zz__zz_S_10) + $signed(_zz__zz_S_10_1));
    _zz_S_11 <= ($signed(_zz__zz_S_11) + $signed(_zz__zz_S_11_1));
    a1Temp_8_regNext <= a1Temp_8;
    _zz_S_12 <= ($signed(_zz__zz_S_12) + $signed(_zz__zz_S_12_1));
    _zz_S_13 <= ($signed(_zz__zz_S_13) + $signed(_zz__zz_S_13_1));
    a1Temp_8_regNext_regNext <= a1Temp_8_regNext;
    _zz_S_14 <= ($signed(_zz__zz_S_14) + $signed(_zz__zz_S_14_1));
    a1Temp_8_regNext_regNext_regNext <= a1Temp_8_regNext_regNext;
    _zz_S_15 <= ($signed(_zz__zz_S_15) + $signed(_zz__zz_S_15_1));
  end


endmodule

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

//WaXpmSyncFifo_1 replaced by WaXpmSyncFifo_1

module WaXpmSyncFifo_1 (
  input               reset,
  input               clk,
  input               dataIn_valid,
  input      [127:0]  dataIn_payload,
  input               rd_en,
  output     [127:0]  dout,
  input               softReset
);

  wire       [127:0]  fifo_dout;
  reg                 dataIn_valid_regNext;
  reg        [127:0]  dataIn_payload_regNext;

  FifoSync_1 fifo (
    .wr_en (dataIn_valid_regNext         ), //i
    .din   (dataIn_payload_regNext[127:0]), //i
    .dout  (fifo_dout[127:0]             ), //o
    .rd_en (rd_en                        ), //i
    .reset (reset                        ), //i
    .clk   (clk                          )  //i
  );
  assign dout = fifo_dout;
  always @(posedge clk) begin
    dataIn_valid_regNext <= dataIn_valid;
    dataIn_payload_regNext <= dataIn_payload;
  end


endmodule

module WaXpmSyncFifo (
  input      [13:0]   sCount,
  input      [13:0]   mCount,
  output reg          sReady,
  output reg          mReady,
  input               reset,
  input               clk,
  input               dataIn_valid,
  input      [127:0]  dataIn_payload,
  input               rd_en,
  output     [127:0]  dout,
  input               softReset
);

  wire       [127:0]  fifo_dout;
  wire       [13:0]   fifo_wr_data_count;
  wire       [13:0]   fifo_rd_data_count;
  wire       [13:0]   _zz_when_WaFifo_l66;
  reg                 dataIn_valid_regNext;
  reg        [127:0]  dataIn_payload_regNext;
  wire                when_WaFifo_l66;
  wire                when_WaFifo_l71;

  assign _zz_when_WaFifo_l66 = (fifo_wr_data_count + sCount);
  FifoSync fifo (
    .wr_en         (dataIn_valid_regNext         ), //i
    .din           (dataIn_payload_regNext[127:0]), //i
    .dout          (fifo_dout[127:0]             ), //o
    .rd_en         (rd_en                        ), //i
    .wr_data_count (fifo_wr_data_count[13:0]     ), //o
    .rd_data_count (fifo_rd_data_count[13:0]     ), //o
    .reset         (reset                        ), //i
    .clk           (clk                          )  //i
  );
  assign dout = fifo_dout;
  assign when_WaFifo_l66 = (_zz_when_WaFifo_l66 < 14'h1ff6);
  assign when_WaFifo_l71 = (mCount <= fifo_rd_data_count);
  always @(posedge clk) begin
    dataIn_valid_regNext <= dataIn_valid;
    dataIn_payload_regNext <= dataIn_payload;
    if(when_WaFifo_l66) begin
      sReady <= 1'b1;
    end else begin
      sReady <= 1'b0;
    end
    if(when_WaFifo_l71) begin
      mReady <= 1'b1;
    end else begin
      mReady <= 1'b0;
    end
  end


endmodule

module LoadWeight (
  input               start,
  input               sData_valid,
  output reg          sData_ready,
  input      [127:0]  sData_payload,
  input      [12:0]   weightNum,
  input      [7:0]    quanNum,
  input      [8:0]    weightRead_0_addr,
  output     [2047:0] weightRead_0_data,
  input      [8:0]    weightRead_1_addr,
  output     [2047:0] weightRead_1_data,
  input      [8:0]    weightRead_2_addr,
  output     [2047:0] weightRead_2_data,
  input      [8:0]    weightRead_3_addr,
  output     [2047:0] weightRead_3_data,
  input      [8:0]    weightRead_4_addr,
  output     [2047:0] weightRead_4_data,
  input      [8:0]    weightRead_5_addr,
  output     [2047:0] weightRead_5_data,
  input      [8:0]    weightRead_6_addr,
  output     [2047:0] weightRead_6_data,
  input      [8:0]    weightRead_7_addr,
  output     [2047:0] weightRead_7_data,
  input      [8:0]    weightRead_8_addr,
  output     [2047:0] weightRead_8_data,
  input      [5:0]    biasRead_addr,
  output     [511:0]  biasRead_data,
  input      [5:0]    scaleRead_addr,
  output     [511:0]  scaleRead_data,
  input      [5:0]    shiftRead_addr,
  output     [511:0]  shiftRead_data,
  output reg          copyWeightDone,
  input      [1:0]    convType,
  input      [11:0]   channelIn,
  input      [11:0]   channelOut,
  input               clk,
  input               reset,
  input               softReset
);
  localparam LoadWeightEnum_IDLE = 6'd1;
  localparam LoadWeightEnum_INIT = 6'd2;
  localparam LoadWeightEnum_COPY_WEIGHT = 6'd4;
  localparam LoadWeightEnum_COPY_BIAS = 6'd8;
  localparam LoadWeightEnum_COPY_SCALE = 6'd16;
  localparam LoadWeightEnum_COPY_SHIFT = 6'd32;

  wire       [8:0]    weightRam_0_0_addra;
  wire       [8:0]    weightRam_0_0_addrb;
  wire       [127:0]  weightRam_0_0_dina;
  wire       [0:0]    weightRam_0_0_wea;
  wire       [8:0]    weightRam_0_1_addra;
  wire       [8:0]    weightRam_0_1_addrb;
  wire       [127:0]  weightRam_0_1_dina;
  wire       [0:0]    weightRam_0_1_wea;
  wire       [8:0]    weightRam_0_2_addra;
  wire       [8:0]    weightRam_0_2_addrb;
  wire       [127:0]  weightRam_0_2_dina;
  wire       [0:0]    weightRam_0_2_wea;
  wire       [8:0]    weightRam_0_3_addra;
  wire       [8:0]    weightRam_0_3_addrb;
  wire       [127:0]  weightRam_0_3_dina;
  wire       [0:0]    weightRam_0_3_wea;
  wire       [8:0]    weightRam_0_4_addra;
  wire       [8:0]    weightRam_0_4_addrb;
  wire       [127:0]  weightRam_0_4_dina;
  wire       [0:0]    weightRam_0_4_wea;
  wire       [8:0]    weightRam_0_5_addra;
  wire       [8:0]    weightRam_0_5_addrb;
  wire       [127:0]  weightRam_0_5_dina;
  wire       [0:0]    weightRam_0_5_wea;
  wire       [8:0]    weightRam_0_6_addra;
  wire       [8:0]    weightRam_0_6_addrb;
  wire       [127:0]  weightRam_0_6_dina;
  wire       [0:0]    weightRam_0_6_wea;
  wire       [8:0]    weightRam_0_7_addra;
  wire       [8:0]    weightRam_0_7_addrb;
  wire       [127:0]  weightRam_0_7_dina;
  wire       [0:0]    weightRam_0_7_wea;
  wire       [8:0]    weightRam_0_8_addra;
  wire       [8:0]    weightRam_0_8_addrb;
  wire       [127:0]  weightRam_0_8_dina;
  wire       [0:0]    weightRam_0_8_wea;
  wire       [8:0]    weightRam_0_9_addra;
  wire       [8:0]    weightRam_0_9_addrb;
  wire       [127:0]  weightRam_0_9_dina;
  wire       [0:0]    weightRam_0_9_wea;
  wire       [8:0]    weightRam_0_10_addra;
  wire       [8:0]    weightRam_0_10_addrb;
  wire       [127:0]  weightRam_0_10_dina;
  wire       [0:0]    weightRam_0_10_wea;
  wire       [8:0]    weightRam_0_11_addra;
  wire       [8:0]    weightRam_0_11_addrb;
  wire       [127:0]  weightRam_0_11_dina;
  wire       [0:0]    weightRam_0_11_wea;
  wire       [8:0]    weightRam_0_12_addra;
  wire       [8:0]    weightRam_0_12_addrb;
  wire       [127:0]  weightRam_0_12_dina;
  wire       [0:0]    weightRam_0_12_wea;
  wire       [8:0]    weightRam_0_13_addra;
  wire       [8:0]    weightRam_0_13_addrb;
  wire       [127:0]  weightRam_0_13_dina;
  wire       [0:0]    weightRam_0_13_wea;
  wire       [8:0]    weightRam_0_14_addra;
  wire       [8:0]    weightRam_0_14_addrb;
  wire       [127:0]  weightRam_0_14_dina;
  wire       [0:0]    weightRam_0_14_wea;
  wire       [8:0]    weightRam_0_15_addra;
  wire       [8:0]    weightRam_0_15_addrb;
  wire       [127:0]  weightRam_0_15_dina;
  wire       [0:0]    weightRam_0_15_wea;
  wire       [8:0]    weightRam_1_0_addra;
  wire       [8:0]    weightRam_1_0_addrb;
  wire       [127:0]  weightRam_1_0_dina;
  wire       [0:0]    weightRam_1_0_wea;
  wire       [8:0]    weightRam_1_1_addra;
  wire       [8:0]    weightRam_1_1_addrb;
  wire       [127:0]  weightRam_1_1_dina;
  wire       [0:0]    weightRam_1_1_wea;
  wire       [8:0]    weightRam_1_2_addra;
  wire       [8:0]    weightRam_1_2_addrb;
  wire       [127:0]  weightRam_1_2_dina;
  wire       [0:0]    weightRam_1_2_wea;
  wire       [8:0]    weightRam_1_3_addra;
  wire       [8:0]    weightRam_1_3_addrb;
  wire       [127:0]  weightRam_1_3_dina;
  wire       [0:0]    weightRam_1_3_wea;
  wire       [8:0]    weightRam_1_4_addra;
  wire       [8:0]    weightRam_1_4_addrb;
  wire       [127:0]  weightRam_1_4_dina;
  wire       [0:0]    weightRam_1_4_wea;
  wire       [8:0]    weightRam_1_5_addra;
  wire       [8:0]    weightRam_1_5_addrb;
  wire       [127:0]  weightRam_1_5_dina;
  wire       [0:0]    weightRam_1_5_wea;
  wire       [8:0]    weightRam_1_6_addra;
  wire       [8:0]    weightRam_1_6_addrb;
  wire       [127:0]  weightRam_1_6_dina;
  wire       [0:0]    weightRam_1_6_wea;
  wire       [8:0]    weightRam_1_7_addra;
  wire       [8:0]    weightRam_1_7_addrb;
  wire       [127:0]  weightRam_1_7_dina;
  wire       [0:0]    weightRam_1_7_wea;
  wire       [8:0]    weightRam_1_8_addra;
  wire       [8:0]    weightRam_1_8_addrb;
  wire       [127:0]  weightRam_1_8_dina;
  wire       [0:0]    weightRam_1_8_wea;
  wire       [8:0]    weightRam_1_9_addra;
  wire       [8:0]    weightRam_1_9_addrb;
  wire       [127:0]  weightRam_1_9_dina;
  wire       [0:0]    weightRam_1_9_wea;
  wire       [8:0]    weightRam_1_10_addra;
  wire       [8:0]    weightRam_1_10_addrb;
  wire       [127:0]  weightRam_1_10_dina;
  wire       [0:0]    weightRam_1_10_wea;
  wire       [8:0]    weightRam_1_11_addra;
  wire       [8:0]    weightRam_1_11_addrb;
  wire       [127:0]  weightRam_1_11_dina;
  wire       [0:0]    weightRam_1_11_wea;
  wire       [8:0]    weightRam_1_12_addra;
  wire       [8:0]    weightRam_1_12_addrb;
  wire       [127:0]  weightRam_1_12_dina;
  wire       [0:0]    weightRam_1_12_wea;
  wire       [8:0]    weightRam_1_13_addra;
  wire       [8:0]    weightRam_1_13_addrb;
  wire       [127:0]  weightRam_1_13_dina;
  wire       [0:0]    weightRam_1_13_wea;
  wire       [8:0]    weightRam_1_14_addra;
  wire       [8:0]    weightRam_1_14_addrb;
  wire       [127:0]  weightRam_1_14_dina;
  wire       [0:0]    weightRam_1_14_wea;
  wire       [8:0]    weightRam_1_15_addra;
  wire       [8:0]    weightRam_1_15_addrb;
  wire       [127:0]  weightRam_1_15_dina;
  wire       [0:0]    weightRam_1_15_wea;
  wire       [8:0]    weightRam_2_0_addra;
  wire       [8:0]    weightRam_2_0_addrb;
  wire       [127:0]  weightRam_2_0_dina;
  wire       [0:0]    weightRam_2_0_wea;
  wire       [8:0]    weightRam_2_1_addra;
  wire       [8:0]    weightRam_2_1_addrb;
  wire       [127:0]  weightRam_2_1_dina;
  wire       [0:0]    weightRam_2_1_wea;
  wire       [8:0]    weightRam_2_2_addra;
  wire       [8:0]    weightRam_2_2_addrb;
  wire       [127:0]  weightRam_2_2_dina;
  wire       [0:0]    weightRam_2_2_wea;
  wire       [8:0]    weightRam_2_3_addra;
  wire       [8:0]    weightRam_2_3_addrb;
  wire       [127:0]  weightRam_2_3_dina;
  wire       [0:0]    weightRam_2_3_wea;
  wire       [8:0]    weightRam_2_4_addra;
  wire       [8:0]    weightRam_2_4_addrb;
  wire       [127:0]  weightRam_2_4_dina;
  wire       [0:0]    weightRam_2_4_wea;
  wire       [8:0]    weightRam_2_5_addra;
  wire       [8:0]    weightRam_2_5_addrb;
  wire       [127:0]  weightRam_2_5_dina;
  wire       [0:0]    weightRam_2_5_wea;
  wire       [8:0]    weightRam_2_6_addra;
  wire       [8:0]    weightRam_2_6_addrb;
  wire       [127:0]  weightRam_2_6_dina;
  wire       [0:0]    weightRam_2_6_wea;
  wire       [8:0]    weightRam_2_7_addra;
  wire       [8:0]    weightRam_2_7_addrb;
  wire       [127:0]  weightRam_2_7_dina;
  wire       [0:0]    weightRam_2_7_wea;
  wire       [8:0]    weightRam_2_8_addra;
  wire       [8:0]    weightRam_2_8_addrb;
  wire       [127:0]  weightRam_2_8_dina;
  wire       [0:0]    weightRam_2_8_wea;
  wire       [8:0]    weightRam_2_9_addra;
  wire       [8:0]    weightRam_2_9_addrb;
  wire       [127:0]  weightRam_2_9_dina;
  wire       [0:0]    weightRam_2_9_wea;
  wire       [8:0]    weightRam_2_10_addra;
  wire       [8:0]    weightRam_2_10_addrb;
  wire       [127:0]  weightRam_2_10_dina;
  wire       [0:0]    weightRam_2_10_wea;
  wire       [8:0]    weightRam_2_11_addra;
  wire       [8:0]    weightRam_2_11_addrb;
  wire       [127:0]  weightRam_2_11_dina;
  wire       [0:0]    weightRam_2_11_wea;
  wire       [8:0]    weightRam_2_12_addra;
  wire       [8:0]    weightRam_2_12_addrb;
  wire       [127:0]  weightRam_2_12_dina;
  wire       [0:0]    weightRam_2_12_wea;
  wire       [8:0]    weightRam_2_13_addra;
  wire       [8:0]    weightRam_2_13_addrb;
  wire       [127:0]  weightRam_2_13_dina;
  wire       [0:0]    weightRam_2_13_wea;
  wire       [8:0]    weightRam_2_14_addra;
  wire       [8:0]    weightRam_2_14_addrb;
  wire       [127:0]  weightRam_2_14_dina;
  wire       [0:0]    weightRam_2_14_wea;
  wire       [8:0]    weightRam_2_15_addra;
  wire       [8:0]    weightRam_2_15_addrb;
  wire       [127:0]  weightRam_2_15_dina;
  wire       [0:0]    weightRam_2_15_wea;
  wire       [8:0]    weightRam_3_0_addra;
  wire       [8:0]    weightRam_3_0_addrb;
  wire       [127:0]  weightRam_3_0_dina;
  wire       [0:0]    weightRam_3_0_wea;
  wire       [8:0]    weightRam_3_1_addra;
  wire       [8:0]    weightRam_3_1_addrb;
  wire       [127:0]  weightRam_3_1_dina;
  wire       [0:0]    weightRam_3_1_wea;
  wire       [8:0]    weightRam_3_2_addra;
  wire       [8:0]    weightRam_3_2_addrb;
  wire       [127:0]  weightRam_3_2_dina;
  wire       [0:0]    weightRam_3_2_wea;
  wire       [8:0]    weightRam_3_3_addra;
  wire       [8:0]    weightRam_3_3_addrb;
  wire       [127:0]  weightRam_3_3_dina;
  wire       [0:0]    weightRam_3_3_wea;
  wire       [8:0]    weightRam_3_4_addra;
  wire       [8:0]    weightRam_3_4_addrb;
  wire       [127:0]  weightRam_3_4_dina;
  wire       [0:0]    weightRam_3_4_wea;
  wire       [8:0]    weightRam_3_5_addra;
  wire       [8:0]    weightRam_3_5_addrb;
  wire       [127:0]  weightRam_3_5_dina;
  wire       [0:0]    weightRam_3_5_wea;
  wire       [8:0]    weightRam_3_6_addra;
  wire       [8:0]    weightRam_3_6_addrb;
  wire       [127:0]  weightRam_3_6_dina;
  wire       [0:0]    weightRam_3_6_wea;
  wire       [8:0]    weightRam_3_7_addra;
  wire       [8:0]    weightRam_3_7_addrb;
  wire       [127:0]  weightRam_3_7_dina;
  wire       [0:0]    weightRam_3_7_wea;
  wire       [8:0]    weightRam_3_8_addra;
  wire       [8:0]    weightRam_3_8_addrb;
  wire       [127:0]  weightRam_3_8_dina;
  wire       [0:0]    weightRam_3_8_wea;
  wire       [8:0]    weightRam_3_9_addra;
  wire       [8:0]    weightRam_3_9_addrb;
  wire       [127:0]  weightRam_3_9_dina;
  wire       [0:0]    weightRam_3_9_wea;
  wire       [8:0]    weightRam_3_10_addra;
  wire       [8:0]    weightRam_3_10_addrb;
  wire       [127:0]  weightRam_3_10_dina;
  wire       [0:0]    weightRam_3_10_wea;
  wire       [8:0]    weightRam_3_11_addra;
  wire       [8:0]    weightRam_3_11_addrb;
  wire       [127:0]  weightRam_3_11_dina;
  wire       [0:0]    weightRam_3_11_wea;
  wire       [8:0]    weightRam_3_12_addra;
  wire       [8:0]    weightRam_3_12_addrb;
  wire       [127:0]  weightRam_3_12_dina;
  wire       [0:0]    weightRam_3_12_wea;
  wire       [8:0]    weightRam_3_13_addra;
  wire       [8:0]    weightRam_3_13_addrb;
  wire       [127:0]  weightRam_3_13_dina;
  wire       [0:0]    weightRam_3_13_wea;
  wire       [8:0]    weightRam_3_14_addra;
  wire       [8:0]    weightRam_3_14_addrb;
  wire       [127:0]  weightRam_3_14_dina;
  wire       [0:0]    weightRam_3_14_wea;
  wire       [8:0]    weightRam_3_15_addra;
  wire       [8:0]    weightRam_3_15_addrb;
  wire       [127:0]  weightRam_3_15_dina;
  wire       [0:0]    weightRam_3_15_wea;
  wire       [8:0]    weightRam_4_0_addra;
  wire       [8:0]    weightRam_4_0_addrb;
  wire       [127:0]  weightRam_4_0_dina;
  wire       [0:0]    weightRam_4_0_wea;
  wire       [8:0]    weightRam_4_1_addra;
  wire       [8:0]    weightRam_4_1_addrb;
  wire       [127:0]  weightRam_4_1_dina;
  wire       [0:0]    weightRam_4_1_wea;
  wire       [8:0]    weightRam_4_2_addra;
  wire       [8:0]    weightRam_4_2_addrb;
  wire       [127:0]  weightRam_4_2_dina;
  wire       [0:0]    weightRam_4_2_wea;
  wire       [8:0]    weightRam_4_3_addra;
  wire       [8:0]    weightRam_4_3_addrb;
  wire       [127:0]  weightRam_4_3_dina;
  wire       [0:0]    weightRam_4_3_wea;
  wire       [8:0]    weightRam_4_4_addra;
  wire       [8:0]    weightRam_4_4_addrb;
  wire       [127:0]  weightRam_4_4_dina;
  wire       [0:0]    weightRam_4_4_wea;
  wire       [8:0]    weightRam_4_5_addra;
  wire       [8:0]    weightRam_4_5_addrb;
  wire       [127:0]  weightRam_4_5_dina;
  wire       [0:0]    weightRam_4_5_wea;
  wire       [8:0]    weightRam_4_6_addra;
  wire       [8:0]    weightRam_4_6_addrb;
  wire       [127:0]  weightRam_4_6_dina;
  wire       [0:0]    weightRam_4_6_wea;
  wire       [8:0]    weightRam_4_7_addra;
  wire       [8:0]    weightRam_4_7_addrb;
  wire       [127:0]  weightRam_4_7_dina;
  wire       [0:0]    weightRam_4_7_wea;
  wire       [8:0]    weightRam_4_8_addra;
  wire       [8:0]    weightRam_4_8_addrb;
  wire       [127:0]  weightRam_4_8_dina;
  wire       [0:0]    weightRam_4_8_wea;
  wire       [8:0]    weightRam_4_9_addra;
  wire       [8:0]    weightRam_4_9_addrb;
  wire       [127:0]  weightRam_4_9_dina;
  wire       [0:0]    weightRam_4_9_wea;
  wire       [8:0]    weightRam_4_10_addra;
  wire       [8:0]    weightRam_4_10_addrb;
  wire       [127:0]  weightRam_4_10_dina;
  wire       [0:0]    weightRam_4_10_wea;
  wire       [8:0]    weightRam_4_11_addra;
  wire       [8:0]    weightRam_4_11_addrb;
  wire       [127:0]  weightRam_4_11_dina;
  wire       [0:0]    weightRam_4_11_wea;
  wire       [8:0]    weightRam_4_12_addra;
  wire       [8:0]    weightRam_4_12_addrb;
  wire       [127:0]  weightRam_4_12_dina;
  wire       [0:0]    weightRam_4_12_wea;
  wire       [8:0]    weightRam_4_13_addra;
  wire       [8:0]    weightRam_4_13_addrb;
  wire       [127:0]  weightRam_4_13_dina;
  wire       [0:0]    weightRam_4_13_wea;
  wire       [8:0]    weightRam_4_14_addra;
  wire       [8:0]    weightRam_4_14_addrb;
  wire       [127:0]  weightRam_4_14_dina;
  wire       [0:0]    weightRam_4_14_wea;
  wire       [8:0]    weightRam_4_15_addra;
  wire       [8:0]    weightRam_4_15_addrb;
  wire       [127:0]  weightRam_4_15_dina;
  wire       [0:0]    weightRam_4_15_wea;
  wire       [8:0]    weightRam_5_0_addra;
  wire       [8:0]    weightRam_5_0_addrb;
  wire       [127:0]  weightRam_5_0_dina;
  wire       [0:0]    weightRam_5_0_wea;
  wire       [8:0]    weightRam_5_1_addra;
  wire       [8:0]    weightRam_5_1_addrb;
  wire       [127:0]  weightRam_5_1_dina;
  wire       [0:0]    weightRam_5_1_wea;
  wire       [8:0]    weightRam_5_2_addra;
  wire       [8:0]    weightRam_5_2_addrb;
  wire       [127:0]  weightRam_5_2_dina;
  wire       [0:0]    weightRam_5_2_wea;
  wire       [8:0]    weightRam_5_3_addra;
  wire       [8:0]    weightRam_5_3_addrb;
  wire       [127:0]  weightRam_5_3_dina;
  wire       [0:0]    weightRam_5_3_wea;
  wire       [8:0]    weightRam_5_4_addra;
  wire       [8:0]    weightRam_5_4_addrb;
  wire       [127:0]  weightRam_5_4_dina;
  wire       [0:0]    weightRam_5_4_wea;
  wire       [8:0]    weightRam_5_5_addra;
  wire       [8:0]    weightRam_5_5_addrb;
  wire       [127:0]  weightRam_5_5_dina;
  wire       [0:0]    weightRam_5_5_wea;
  wire       [8:0]    weightRam_5_6_addra;
  wire       [8:0]    weightRam_5_6_addrb;
  wire       [127:0]  weightRam_5_6_dina;
  wire       [0:0]    weightRam_5_6_wea;
  wire       [8:0]    weightRam_5_7_addra;
  wire       [8:0]    weightRam_5_7_addrb;
  wire       [127:0]  weightRam_5_7_dina;
  wire       [0:0]    weightRam_5_7_wea;
  wire       [8:0]    weightRam_5_8_addra;
  wire       [8:0]    weightRam_5_8_addrb;
  wire       [127:0]  weightRam_5_8_dina;
  wire       [0:0]    weightRam_5_8_wea;
  wire       [8:0]    weightRam_5_9_addra;
  wire       [8:0]    weightRam_5_9_addrb;
  wire       [127:0]  weightRam_5_9_dina;
  wire       [0:0]    weightRam_5_9_wea;
  wire       [8:0]    weightRam_5_10_addra;
  wire       [8:0]    weightRam_5_10_addrb;
  wire       [127:0]  weightRam_5_10_dina;
  wire       [0:0]    weightRam_5_10_wea;
  wire       [8:0]    weightRam_5_11_addra;
  wire       [8:0]    weightRam_5_11_addrb;
  wire       [127:0]  weightRam_5_11_dina;
  wire       [0:0]    weightRam_5_11_wea;
  wire       [8:0]    weightRam_5_12_addra;
  wire       [8:0]    weightRam_5_12_addrb;
  wire       [127:0]  weightRam_5_12_dina;
  wire       [0:0]    weightRam_5_12_wea;
  wire       [8:0]    weightRam_5_13_addra;
  wire       [8:0]    weightRam_5_13_addrb;
  wire       [127:0]  weightRam_5_13_dina;
  wire       [0:0]    weightRam_5_13_wea;
  wire       [8:0]    weightRam_5_14_addra;
  wire       [8:0]    weightRam_5_14_addrb;
  wire       [127:0]  weightRam_5_14_dina;
  wire       [0:0]    weightRam_5_14_wea;
  wire       [8:0]    weightRam_5_15_addra;
  wire       [8:0]    weightRam_5_15_addrb;
  wire       [127:0]  weightRam_5_15_dina;
  wire       [0:0]    weightRam_5_15_wea;
  wire       [8:0]    weightRam_6_0_addra;
  wire       [8:0]    weightRam_6_0_addrb;
  wire       [127:0]  weightRam_6_0_dina;
  wire       [0:0]    weightRam_6_0_wea;
  wire       [8:0]    weightRam_6_1_addra;
  wire       [8:0]    weightRam_6_1_addrb;
  wire       [127:0]  weightRam_6_1_dina;
  wire       [0:0]    weightRam_6_1_wea;
  wire       [8:0]    weightRam_6_2_addra;
  wire       [8:0]    weightRam_6_2_addrb;
  wire       [127:0]  weightRam_6_2_dina;
  wire       [0:0]    weightRam_6_2_wea;
  wire       [8:0]    weightRam_6_3_addra;
  wire       [8:0]    weightRam_6_3_addrb;
  wire       [127:0]  weightRam_6_3_dina;
  wire       [0:0]    weightRam_6_3_wea;
  wire       [8:0]    weightRam_6_4_addra;
  wire       [8:0]    weightRam_6_4_addrb;
  wire       [127:0]  weightRam_6_4_dina;
  wire       [0:0]    weightRam_6_4_wea;
  wire       [8:0]    weightRam_6_5_addra;
  wire       [8:0]    weightRam_6_5_addrb;
  wire       [127:0]  weightRam_6_5_dina;
  wire       [0:0]    weightRam_6_5_wea;
  wire       [8:0]    weightRam_6_6_addra;
  wire       [8:0]    weightRam_6_6_addrb;
  wire       [127:0]  weightRam_6_6_dina;
  wire       [0:0]    weightRam_6_6_wea;
  wire       [8:0]    weightRam_6_7_addra;
  wire       [8:0]    weightRam_6_7_addrb;
  wire       [127:0]  weightRam_6_7_dina;
  wire       [0:0]    weightRam_6_7_wea;
  wire       [8:0]    weightRam_6_8_addra;
  wire       [8:0]    weightRam_6_8_addrb;
  wire       [127:0]  weightRam_6_8_dina;
  wire       [0:0]    weightRam_6_8_wea;
  wire       [8:0]    weightRam_6_9_addra;
  wire       [8:0]    weightRam_6_9_addrb;
  wire       [127:0]  weightRam_6_9_dina;
  wire       [0:0]    weightRam_6_9_wea;
  wire       [8:0]    weightRam_6_10_addra;
  wire       [8:0]    weightRam_6_10_addrb;
  wire       [127:0]  weightRam_6_10_dina;
  wire       [0:0]    weightRam_6_10_wea;
  wire       [8:0]    weightRam_6_11_addra;
  wire       [8:0]    weightRam_6_11_addrb;
  wire       [127:0]  weightRam_6_11_dina;
  wire       [0:0]    weightRam_6_11_wea;
  wire       [8:0]    weightRam_6_12_addra;
  wire       [8:0]    weightRam_6_12_addrb;
  wire       [127:0]  weightRam_6_12_dina;
  wire       [0:0]    weightRam_6_12_wea;
  wire       [8:0]    weightRam_6_13_addra;
  wire       [8:0]    weightRam_6_13_addrb;
  wire       [127:0]  weightRam_6_13_dina;
  wire       [0:0]    weightRam_6_13_wea;
  wire       [8:0]    weightRam_6_14_addra;
  wire       [8:0]    weightRam_6_14_addrb;
  wire       [127:0]  weightRam_6_14_dina;
  wire       [0:0]    weightRam_6_14_wea;
  wire       [8:0]    weightRam_6_15_addra;
  wire       [8:0]    weightRam_6_15_addrb;
  wire       [127:0]  weightRam_6_15_dina;
  wire       [0:0]    weightRam_6_15_wea;
  wire       [8:0]    weightRam_7_0_addra;
  wire       [8:0]    weightRam_7_0_addrb;
  wire       [127:0]  weightRam_7_0_dina;
  wire       [0:0]    weightRam_7_0_wea;
  wire       [8:0]    weightRam_7_1_addra;
  wire       [8:0]    weightRam_7_1_addrb;
  wire       [127:0]  weightRam_7_1_dina;
  wire       [0:0]    weightRam_7_1_wea;
  wire       [8:0]    weightRam_7_2_addra;
  wire       [8:0]    weightRam_7_2_addrb;
  wire       [127:0]  weightRam_7_2_dina;
  wire       [0:0]    weightRam_7_2_wea;
  wire       [8:0]    weightRam_7_3_addra;
  wire       [8:0]    weightRam_7_3_addrb;
  wire       [127:0]  weightRam_7_3_dina;
  wire       [0:0]    weightRam_7_3_wea;
  wire       [8:0]    weightRam_7_4_addra;
  wire       [8:0]    weightRam_7_4_addrb;
  wire       [127:0]  weightRam_7_4_dina;
  wire       [0:0]    weightRam_7_4_wea;
  wire       [8:0]    weightRam_7_5_addra;
  wire       [8:0]    weightRam_7_5_addrb;
  wire       [127:0]  weightRam_7_5_dina;
  wire       [0:0]    weightRam_7_5_wea;
  wire       [8:0]    weightRam_7_6_addra;
  wire       [8:0]    weightRam_7_6_addrb;
  wire       [127:0]  weightRam_7_6_dina;
  wire       [0:0]    weightRam_7_6_wea;
  wire       [8:0]    weightRam_7_7_addra;
  wire       [8:0]    weightRam_7_7_addrb;
  wire       [127:0]  weightRam_7_7_dina;
  wire       [0:0]    weightRam_7_7_wea;
  wire       [8:0]    weightRam_7_8_addra;
  wire       [8:0]    weightRam_7_8_addrb;
  wire       [127:0]  weightRam_7_8_dina;
  wire       [0:0]    weightRam_7_8_wea;
  wire       [8:0]    weightRam_7_9_addra;
  wire       [8:0]    weightRam_7_9_addrb;
  wire       [127:0]  weightRam_7_9_dina;
  wire       [0:0]    weightRam_7_9_wea;
  wire       [8:0]    weightRam_7_10_addra;
  wire       [8:0]    weightRam_7_10_addrb;
  wire       [127:0]  weightRam_7_10_dina;
  wire       [0:0]    weightRam_7_10_wea;
  wire       [8:0]    weightRam_7_11_addra;
  wire       [8:0]    weightRam_7_11_addrb;
  wire       [127:0]  weightRam_7_11_dina;
  wire       [0:0]    weightRam_7_11_wea;
  wire       [8:0]    weightRam_7_12_addra;
  wire       [8:0]    weightRam_7_12_addrb;
  wire       [127:0]  weightRam_7_12_dina;
  wire       [0:0]    weightRam_7_12_wea;
  wire       [8:0]    weightRam_7_13_addra;
  wire       [8:0]    weightRam_7_13_addrb;
  wire       [127:0]  weightRam_7_13_dina;
  wire       [0:0]    weightRam_7_13_wea;
  wire       [8:0]    weightRam_7_14_addra;
  wire       [8:0]    weightRam_7_14_addrb;
  wire       [127:0]  weightRam_7_14_dina;
  wire       [0:0]    weightRam_7_14_wea;
  wire       [8:0]    weightRam_7_15_addra;
  wire       [8:0]    weightRam_7_15_addrb;
  wire       [127:0]  weightRam_7_15_dina;
  wire       [0:0]    weightRam_7_15_wea;
  wire       [8:0]    weightRam_8_0_addra;
  wire       [8:0]    weightRam_8_0_addrb;
  wire       [127:0]  weightRam_8_0_dina;
  wire       [0:0]    weightRam_8_0_wea;
  wire       [8:0]    weightRam_8_1_addra;
  wire       [8:0]    weightRam_8_1_addrb;
  wire       [127:0]  weightRam_8_1_dina;
  wire       [0:0]    weightRam_8_1_wea;
  wire       [8:0]    weightRam_8_2_addra;
  wire       [8:0]    weightRam_8_2_addrb;
  wire       [127:0]  weightRam_8_2_dina;
  wire       [0:0]    weightRam_8_2_wea;
  wire       [8:0]    weightRam_8_3_addra;
  wire       [8:0]    weightRam_8_3_addrb;
  wire       [127:0]  weightRam_8_3_dina;
  wire       [0:0]    weightRam_8_3_wea;
  wire       [8:0]    weightRam_8_4_addra;
  wire       [8:0]    weightRam_8_4_addrb;
  wire       [127:0]  weightRam_8_4_dina;
  wire       [0:0]    weightRam_8_4_wea;
  wire       [8:0]    weightRam_8_5_addra;
  wire       [8:0]    weightRam_8_5_addrb;
  wire       [127:0]  weightRam_8_5_dina;
  wire       [0:0]    weightRam_8_5_wea;
  wire       [8:0]    weightRam_8_6_addra;
  wire       [8:0]    weightRam_8_6_addrb;
  wire       [127:0]  weightRam_8_6_dina;
  wire       [0:0]    weightRam_8_6_wea;
  wire       [8:0]    weightRam_8_7_addra;
  wire       [8:0]    weightRam_8_7_addrb;
  wire       [127:0]  weightRam_8_7_dina;
  wire       [0:0]    weightRam_8_7_wea;
  wire       [8:0]    weightRam_8_8_addra;
  wire       [8:0]    weightRam_8_8_addrb;
  wire       [127:0]  weightRam_8_8_dina;
  wire       [0:0]    weightRam_8_8_wea;
  wire       [8:0]    weightRam_8_9_addra;
  wire       [8:0]    weightRam_8_9_addrb;
  wire       [127:0]  weightRam_8_9_dina;
  wire       [0:0]    weightRam_8_9_wea;
  wire       [8:0]    weightRam_8_10_addra;
  wire       [8:0]    weightRam_8_10_addrb;
  wire       [127:0]  weightRam_8_10_dina;
  wire       [0:0]    weightRam_8_10_wea;
  wire       [8:0]    weightRam_8_11_addra;
  wire       [8:0]    weightRam_8_11_addrb;
  wire       [127:0]  weightRam_8_11_dina;
  wire       [0:0]    weightRam_8_11_wea;
  wire       [8:0]    weightRam_8_12_addra;
  wire       [8:0]    weightRam_8_12_addrb;
  wire       [127:0]  weightRam_8_12_dina;
  wire       [0:0]    weightRam_8_12_wea;
  wire       [8:0]    weightRam_8_13_addra;
  wire       [8:0]    weightRam_8_13_addrb;
  wire       [127:0]  weightRam_8_13_dina;
  wire       [0:0]    weightRam_8_13_wea;
  wire       [8:0]    weightRam_8_14_addra;
  wire       [8:0]    weightRam_8_14_addrb;
  wire       [127:0]  weightRam_8_14_dina;
  wire       [0:0]    weightRam_8_14_wea;
  wire       [8:0]    weightRam_8_15_addra;
  wire       [8:0]    weightRam_8_15_addrb;
  wire       [127:0]  weightRam_8_15_dina;
  wire       [0:0]    weightRam_8_15_wea;
  wire       [7:0]    copyBias_ram_addra;
  wire       [5:0]    copyBias_ram_addrb;
  wire       [127:0]  copyBias_ram_dina;
  wire       [0:0]    copyBias_ram_wea;
  wire       [7:0]    copyScale_ram_addra;
  wire       [5:0]    copyScale_ram_addrb;
  wire       [127:0]  copyScale_ram_dina;
  wire       [0:0]    copyScale_ram_wea;
  wire       [7:0]    copyShift_ram_addra;
  wire       [5:0]    copyShift_ram_addrb;
  wire       [127:0]  copyShift_ram_dina;
  wire       [0:0]    copyShift_ram_wea;
  wire       [127:0]  weightRam_0_0_doutb;
  wire       [127:0]  weightRam_0_1_doutb;
  wire       [127:0]  weightRam_0_2_doutb;
  wire       [127:0]  weightRam_0_3_doutb;
  wire       [127:0]  weightRam_0_4_doutb;
  wire       [127:0]  weightRam_0_5_doutb;
  wire       [127:0]  weightRam_0_6_doutb;
  wire       [127:0]  weightRam_0_7_doutb;
  wire       [127:0]  weightRam_0_8_doutb;
  wire       [127:0]  weightRam_0_9_doutb;
  wire       [127:0]  weightRam_0_10_doutb;
  wire       [127:0]  weightRam_0_11_doutb;
  wire       [127:0]  weightRam_0_12_doutb;
  wire       [127:0]  weightRam_0_13_doutb;
  wire       [127:0]  weightRam_0_14_doutb;
  wire       [127:0]  weightRam_0_15_doutb;
  wire       [127:0]  weightRam_1_0_doutb;
  wire       [127:0]  weightRam_1_1_doutb;
  wire       [127:0]  weightRam_1_2_doutb;
  wire       [127:0]  weightRam_1_3_doutb;
  wire       [127:0]  weightRam_1_4_doutb;
  wire       [127:0]  weightRam_1_5_doutb;
  wire       [127:0]  weightRam_1_6_doutb;
  wire       [127:0]  weightRam_1_7_doutb;
  wire       [127:0]  weightRam_1_8_doutb;
  wire       [127:0]  weightRam_1_9_doutb;
  wire       [127:0]  weightRam_1_10_doutb;
  wire       [127:0]  weightRam_1_11_doutb;
  wire       [127:0]  weightRam_1_12_doutb;
  wire       [127:0]  weightRam_1_13_doutb;
  wire       [127:0]  weightRam_1_14_doutb;
  wire       [127:0]  weightRam_1_15_doutb;
  wire       [127:0]  weightRam_2_0_doutb;
  wire       [127:0]  weightRam_2_1_doutb;
  wire       [127:0]  weightRam_2_2_doutb;
  wire       [127:0]  weightRam_2_3_doutb;
  wire       [127:0]  weightRam_2_4_doutb;
  wire       [127:0]  weightRam_2_5_doutb;
  wire       [127:0]  weightRam_2_6_doutb;
  wire       [127:0]  weightRam_2_7_doutb;
  wire       [127:0]  weightRam_2_8_doutb;
  wire       [127:0]  weightRam_2_9_doutb;
  wire       [127:0]  weightRam_2_10_doutb;
  wire       [127:0]  weightRam_2_11_doutb;
  wire       [127:0]  weightRam_2_12_doutb;
  wire       [127:0]  weightRam_2_13_doutb;
  wire       [127:0]  weightRam_2_14_doutb;
  wire       [127:0]  weightRam_2_15_doutb;
  wire       [127:0]  weightRam_3_0_doutb;
  wire       [127:0]  weightRam_3_1_doutb;
  wire       [127:0]  weightRam_3_2_doutb;
  wire       [127:0]  weightRam_3_3_doutb;
  wire       [127:0]  weightRam_3_4_doutb;
  wire       [127:0]  weightRam_3_5_doutb;
  wire       [127:0]  weightRam_3_6_doutb;
  wire       [127:0]  weightRam_3_7_doutb;
  wire       [127:0]  weightRam_3_8_doutb;
  wire       [127:0]  weightRam_3_9_doutb;
  wire       [127:0]  weightRam_3_10_doutb;
  wire       [127:0]  weightRam_3_11_doutb;
  wire       [127:0]  weightRam_3_12_doutb;
  wire       [127:0]  weightRam_3_13_doutb;
  wire       [127:0]  weightRam_3_14_doutb;
  wire       [127:0]  weightRam_3_15_doutb;
  wire       [127:0]  weightRam_4_0_doutb;
  wire       [127:0]  weightRam_4_1_doutb;
  wire       [127:0]  weightRam_4_2_doutb;
  wire       [127:0]  weightRam_4_3_doutb;
  wire       [127:0]  weightRam_4_4_doutb;
  wire       [127:0]  weightRam_4_5_doutb;
  wire       [127:0]  weightRam_4_6_doutb;
  wire       [127:0]  weightRam_4_7_doutb;
  wire       [127:0]  weightRam_4_8_doutb;
  wire       [127:0]  weightRam_4_9_doutb;
  wire       [127:0]  weightRam_4_10_doutb;
  wire       [127:0]  weightRam_4_11_doutb;
  wire       [127:0]  weightRam_4_12_doutb;
  wire       [127:0]  weightRam_4_13_doutb;
  wire       [127:0]  weightRam_4_14_doutb;
  wire       [127:0]  weightRam_4_15_doutb;
  wire       [127:0]  weightRam_5_0_doutb;
  wire       [127:0]  weightRam_5_1_doutb;
  wire       [127:0]  weightRam_5_2_doutb;
  wire       [127:0]  weightRam_5_3_doutb;
  wire       [127:0]  weightRam_5_4_doutb;
  wire       [127:0]  weightRam_5_5_doutb;
  wire       [127:0]  weightRam_5_6_doutb;
  wire       [127:0]  weightRam_5_7_doutb;
  wire       [127:0]  weightRam_5_8_doutb;
  wire       [127:0]  weightRam_5_9_doutb;
  wire       [127:0]  weightRam_5_10_doutb;
  wire       [127:0]  weightRam_5_11_doutb;
  wire       [127:0]  weightRam_5_12_doutb;
  wire       [127:0]  weightRam_5_13_doutb;
  wire       [127:0]  weightRam_5_14_doutb;
  wire       [127:0]  weightRam_5_15_doutb;
  wire       [127:0]  weightRam_6_0_doutb;
  wire       [127:0]  weightRam_6_1_doutb;
  wire       [127:0]  weightRam_6_2_doutb;
  wire       [127:0]  weightRam_6_3_doutb;
  wire       [127:0]  weightRam_6_4_doutb;
  wire       [127:0]  weightRam_6_5_doutb;
  wire       [127:0]  weightRam_6_6_doutb;
  wire       [127:0]  weightRam_6_7_doutb;
  wire       [127:0]  weightRam_6_8_doutb;
  wire       [127:0]  weightRam_6_9_doutb;
  wire       [127:0]  weightRam_6_10_doutb;
  wire       [127:0]  weightRam_6_11_doutb;
  wire       [127:0]  weightRam_6_12_doutb;
  wire       [127:0]  weightRam_6_13_doutb;
  wire       [127:0]  weightRam_6_14_doutb;
  wire       [127:0]  weightRam_6_15_doutb;
  wire       [127:0]  weightRam_7_0_doutb;
  wire       [127:0]  weightRam_7_1_doutb;
  wire       [127:0]  weightRam_7_2_doutb;
  wire       [127:0]  weightRam_7_3_doutb;
  wire       [127:0]  weightRam_7_4_doutb;
  wire       [127:0]  weightRam_7_5_doutb;
  wire       [127:0]  weightRam_7_6_doutb;
  wire       [127:0]  weightRam_7_7_doutb;
  wire       [127:0]  weightRam_7_8_doutb;
  wire       [127:0]  weightRam_7_9_doutb;
  wire       [127:0]  weightRam_7_10_doutb;
  wire       [127:0]  weightRam_7_11_doutb;
  wire       [127:0]  weightRam_7_12_doutb;
  wire       [127:0]  weightRam_7_13_doutb;
  wire       [127:0]  weightRam_7_14_doutb;
  wire       [127:0]  weightRam_7_15_doutb;
  wire       [127:0]  weightRam_8_0_doutb;
  wire       [127:0]  weightRam_8_1_doutb;
  wire       [127:0]  weightRam_8_2_doutb;
  wire       [127:0]  weightRam_8_3_doutb;
  wire       [127:0]  weightRam_8_4_doutb;
  wire       [127:0]  weightRam_8_5_doutb;
  wire       [127:0]  weightRam_8_6_doutb;
  wire       [127:0]  weightRam_8_7_doutb;
  wire       [127:0]  weightRam_8_8_doutb;
  wire       [127:0]  weightRam_8_9_doutb;
  wire       [127:0]  weightRam_8_10_doutb;
  wire       [127:0]  weightRam_8_11_doutb;
  wire       [127:0]  weightRam_8_12_doutb;
  wire       [127:0]  weightRam_8_13_doutb;
  wire       [127:0]  weightRam_8_14_doutb;
  wire       [127:0]  weightRam_8_15_doutb;
  wire       [511:0]  copyBias_ram_doutb;
  wire       [511:0]  copyScale_ram_doutb;
  wire       [511:0]  copyShift_ram_doutb;
  wire       [12:0]   _zz_when_WaCounter_l12_1;
  wire       [7:0]    _zz_when_WaCounter_l12_3;
  wire       [11:0]   _zz_when_WaCounter_l12_6;
  wire       [12:0]   _zz_when_Weight_l326;
  wire       [12:0]   _zz_when_Weight_l326_1;
  wire       [12:0]   _zz_when_Weight_l326_2;
  wire       [12:0]   _zz_when_Weight_l326_3;
  wire       [12:0]   _zz_when_Weight_l326_4;
  wire       [12:0]   _zz_when_Weight_l326_5;
  wire       [12:0]   _zz_when_Weight_l326_6;
  wire       [12:0]   _zz_when_Weight_l326_7;
  wire       [12:0]   _zz_when_Weight_l326_8;
  wire       [12:0]   _zz_when_Weight_l326_9;
  wire       [12:0]   _zz_when_Weight_l326_10;
  wire       [12:0]   _zz_when_Weight_l326_11;
  wire       [12:0]   _zz_when_Weight_l326_12;
  wire       [12:0]   _zz_when_Weight_l326_13;
  wire       [12:0]   _zz_when_Weight_l326_14;
  wire       [12:0]   _zz_when_Weight_l326_15;
  wire       [12:0]   _zz_when_Weight_l326_16;
  wire       [12:0]   _zz_when_Weight_l326_17;
  wire       [12:0]   _zz_when_Weight_l326_18;
  wire       [12:0]   _zz_when_Weight_l326_19;
  wire       [12:0]   _zz_when_Weight_l326_20;
  wire       [12:0]   _zz_when_Weight_l326_21;
  wire       [12:0]   _zz_when_Weight_l326_22;
  wire       [12:0]   _zz_when_Weight_l326_23;
  wire       [12:0]   _zz_when_Weight_l326_24;
  wire       [12:0]   _zz_when_Weight_l326_25;
  wire       [12:0]   _zz_when_Weight_l326_26;
  wire       [12:0]   _zz_when_Weight_l326_27;
  wire       [12:0]   _zz_when_Weight_l326_28;
  wire       [12:0]   _zz_when_Weight_l326_29;
  wire       [12:0]   _zz_when_Weight_l326_30;
  wire       [12:0]   _zz_when_Weight_l326_31;
  wire       [12:0]   _zz_when_Weight_l326_32;
  wire       [12:0]   _zz_when_Weight_l326_33;
  wire       [12:0]   _zz_when_Weight_l326_34;
  wire       [12:0]   _zz_when_Weight_l326_35;
  wire       [12:0]   _zz_when_Weight_l326_36;
  wire       [12:0]   _zz_when_Weight_l326_37;
  wire       [12:0]   _zz_when_Weight_l326_38;
  wire       [12:0]   _zz_when_Weight_l326_39;
  wire       [12:0]   _zz_when_Weight_l326_40;
  wire       [12:0]   _zz_when_Weight_l326_41;
  wire       [12:0]   _zz_when_Weight_l326_42;
  wire       [12:0]   _zz_when_Weight_l326_43;
  wire       [12:0]   _zz_when_Weight_l326_44;
  wire       [12:0]   _zz_when_Weight_l326_45;
  wire       [12:0]   _zz_when_Weight_l326_46;
  wire       [12:0]   _zz_when_Weight_l326_47;
  wire       [12:0]   _zz_when_Weight_l326_48;
  wire       [12:0]   _zz_when_Weight_l326_49;
  wire       [12:0]   _zz_when_Weight_l326_50;
  wire       [12:0]   _zz_when_Weight_l326_51;
  wire       [12:0]   _zz_when_Weight_l326_52;
  wire       [12:0]   _zz_when_Weight_l326_53;
  wire       [12:0]   _zz_when_Weight_l326_54;
  wire       [12:0]   _zz_when_Weight_l326_55;
  wire       [12:0]   _zz_when_Weight_l326_56;
  wire       [12:0]   _zz_when_Weight_l326_57;
  wire       [12:0]   _zz_when_Weight_l326_58;
  wire       [12:0]   _zz_when_Weight_l326_59;
  wire       [12:0]   _zz_when_Weight_l326_60;
  wire       [12:0]   _zz_when_Weight_l326_61;
  wire       [12:0]   _zz_when_Weight_l326_62;
  wire       [12:0]   _zz_when_Weight_l326_63;
  wire       [12:0]   _zz_when_Weight_l326_64;
  wire       [12:0]   _zz_when_Weight_l326_65;
  wire       [12:0]   _zz_when_Weight_l326_66;
  wire       [12:0]   _zz_when_Weight_l326_67;
  wire       [12:0]   _zz_when_Weight_l326_68;
  wire       [12:0]   _zz_when_Weight_l326_69;
  wire       [12:0]   _zz_when_Weight_l326_70;
  wire       [12:0]   _zz_when_Weight_l326_71;
  wire       [12:0]   _zz_when_Weight_l326_72;
  wire       [12:0]   _zz_when_Weight_l326_73;
  wire       [12:0]   _zz_when_Weight_l326_74;
  wire       [12:0]   _zz_when_Weight_l326_75;
  wire       [12:0]   _zz_when_Weight_l326_76;
  wire       [12:0]   _zz_when_Weight_l326_77;
  wire       [12:0]   _zz_when_Weight_l326_78;
  wire       [12:0]   _zz_when_Weight_l326_79;
  wire       [12:0]   _zz_when_Weight_l326_80;
  wire       [12:0]   _zz_when_Weight_l326_81;
  wire       [12:0]   _zz_when_Weight_l326_82;
  wire       [12:0]   _zz_when_Weight_l326_83;
  wire       [12:0]   _zz_when_Weight_l326_84;
  wire       [12:0]   _zz_when_Weight_l326_85;
  wire       [12:0]   _zz_when_Weight_l326_86;
  wire       [12:0]   _zz_when_Weight_l326_87;
  wire       [12:0]   _zz_when_Weight_l326_88;
  wire       [12:0]   _zz_when_Weight_l326_89;
  wire       [12:0]   _zz_when_Weight_l326_90;
  wire       [12:0]   _zz_when_Weight_l326_91;
  wire       [12:0]   _zz_when_Weight_l326_92;
  wire       [12:0]   _zz_when_Weight_l326_93;
  wire       [12:0]   _zz_when_Weight_l326_94;
  wire       [12:0]   _zz_when_Weight_l326_95;
  wire       [12:0]   _zz_when_Weight_l326_96;
  wire       [12:0]   _zz_when_Weight_l326_97;
  wire       [12:0]   _zz_when_Weight_l326_98;
  wire       [12:0]   _zz_when_Weight_l326_99;
  wire       [12:0]   _zz_when_Weight_l326_100;
  wire       [12:0]   _zz_when_Weight_l326_101;
  wire       [12:0]   _zz_when_Weight_l326_102;
  wire       [12:0]   _zz_when_Weight_l326_103;
  wire       [12:0]   _zz_when_Weight_l326_104;
  wire       [12:0]   _zz_when_Weight_l326_105;
  wire       [12:0]   _zz_when_Weight_l326_106;
  wire       [12:0]   _zz_when_Weight_l326_107;
  wire       [12:0]   _zz_when_Weight_l326_108;
  wire       [12:0]   _zz_when_Weight_l326_109;
  wire       [12:0]   _zz_when_Weight_l326_110;
  wire       [12:0]   _zz_when_Weight_l326_111;
  wire       [12:0]   _zz_when_Weight_l326_112;
  wire       [12:0]   _zz_when_Weight_l326_113;
  wire       [12:0]   _zz_when_Weight_l326_114;
  wire       [12:0]   _zz_when_Weight_l326_115;
  wire       [12:0]   _zz_when_Weight_l326_116;
  wire       [12:0]   _zz_when_Weight_l326_117;
  wire       [12:0]   _zz_when_Weight_l326_118;
  wire       [12:0]   _zz_when_Weight_l326_119;
  wire       [12:0]   _zz_when_Weight_l326_120;
  wire       [12:0]   _zz_when_Weight_l326_121;
  wire       [12:0]   _zz_when_Weight_l326_122;
  wire       [12:0]   _zz_when_Weight_l326_123;
  wire       [12:0]   _zz_when_Weight_l326_124;
  wire       [12:0]   _zz_when_Weight_l326_125;
  wire       [12:0]   _zz_when_Weight_l326_126;
  wire       [12:0]   _zz_when_Weight_l326_127;
  wire       [12:0]   _zz_when_Weight_l326_128;
  wire       [12:0]   _zz_when_Weight_l326_129;
  wire       [12:0]   _zz_when_Weight_l326_130;
  wire       [12:0]   _zz_when_Weight_l326_131;
  wire       [12:0]   _zz_when_Weight_l326_132;
  wire       [12:0]   _zz_when_Weight_l326_133;
  wire       [12:0]   _zz_when_Weight_l326_134;
  wire       [12:0]   _zz_when_Weight_l326_135;
  wire       [12:0]   _zz_when_Weight_l326_136;
  wire       [12:0]   _zz_when_Weight_l326_137;
  wire       [12:0]   _zz_when_Weight_l326_138;
  wire       [12:0]   _zz_when_Weight_l326_139;
  wire       [12:0]   _zz_when_Weight_l326_140;
  wire       [12:0]   _zz_when_Weight_l326_141;
  wire       [12:0]   _zz_when_Weight_l326_142;
  wire       [12:0]   _zz_when_Weight_l326_143;
  wire       [1279:0] _zz_weightRead_0_data;
  wire       [383:0]  _zz_weightRead_0_data_1;
  wire       [127:0]  _zz_weightRead_0_data_2;
  wire       [1279:0] _zz_weightRead_1_data;
  wire       [383:0]  _zz_weightRead_1_data_1;
  wire       [127:0]  _zz_weightRead_1_data_2;
  wire       [1279:0] _zz_weightRead_2_data;
  wire       [383:0]  _zz_weightRead_2_data_1;
  wire       [127:0]  _zz_weightRead_2_data_2;
  wire       [1279:0] _zz_weightRead_3_data;
  wire       [383:0]  _zz_weightRead_3_data_1;
  wire       [127:0]  _zz_weightRead_3_data_2;
  wire       [1279:0] _zz_weightRead_4_data;
  wire       [383:0]  _zz_weightRead_4_data_1;
  wire       [127:0]  _zz_weightRead_4_data_2;
  wire       [1279:0] _zz_weightRead_5_data;
  wire       [383:0]  _zz_weightRead_5_data_1;
  wire       [127:0]  _zz_weightRead_5_data_2;
  wire       [1279:0] _zz_weightRead_6_data;
  wire       [383:0]  _zz_weightRead_6_data_1;
  wire       [127:0]  _zz_weightRead_6_data_2;
  wire       [1279:0] _zz_weightRead_7_data;
  wire       [383:0]  _zz_weightRead_7_data_1;
  wire       [127:0]  _zz_weightRead_7_data_2;
  wire       [1279:0] _zz_weightRead_8_data;
  wire       [383:0]  _zz_weightRead_8_data_1;
  wire       [127:0]  _zz_weightRead_8_data_2;
  wire       [12:0]   _zz_addra;
  wire       [12:0]   _zz_addra_1;
  wire       [12:0]   _zz_addra_2;
  wire       [12:0]   _zz_addra_3;
  wire       [12:0]   _zz_addra_4;
  wire       [12:0]   _zz_addra_5;
  wire       [12:0]   _zz_addra_6;
  wire       [12:0]   _zz_addra_7;
  wire       [12:0]   _zz_addra_8;
  wire       [12:0]   _zz_addra_9;
  wire       [12:0]   _zz_addra_10;
  wire       [12:0]   _zz_addra_11;
  wire       [12:0]   _zz_addra_12;
  wire       [12:0]   _zz_addra_13;
  wire       [12:0]   _zz_addra_14;
  wire       [12:0]   _zz_addra_15;
  wire       [12:0]   _zz_addra_16;
  wire       [12:0]   _zz_addra_17;
  wire       [12:0]   _zz_addra_18;
  wire       [12:0]   _zz_addra_19;
  wire       [12:0]   _zz_addra_20;
  wire       [12:0]   _zz_addra_21;
  wire       [12:0]   _zz_addra_22;
  wire       [12:0]   _zz_addra_23;
  wire       [12:0]   _zz_addra_24;
  wire       [12:0]   _zz_addra_25;
  wire       [12:0]   _zz_addra_26;
  wire       [12:0]   _zz_addra_27;
  wire       [12:0]   _zz_addra_28;
  wire       [12:0]   _zz_addra_29;
  wire       [12:0]   _zz_addra_30;
  wire       [12:0]   _zz_addra_31;
  wire       [12:0]   _zz_addra_32;
  wire       [12:0]   _zz_addra_33;
  wire       [12:0]   _zz_addra_34;
  wire       [12:0]   _zz_addra_35;
  wire       [12:0]   _zz_addra_36;
  wire       [12:0]   _zz_addra_37;
  wire       [12:0]   _zz_addra_38;
  wire       [12:0]   _zz_addra_39;
  wire       [12:0]   _zz_addra_40;
  wire       [12:0]   _zz_addra_41;
  wire       [12:0]   _zz_addra_42;
  wire       [12:0]   _zz_addra_43;
  wire       [12:0]   _zz_addra_44;
  wire       [12:0]   _zz_addra_45;
  wire       [12:0]   _zz_addra_46;
  wire       [12:0]   _zz_addra_47;
  wire       [12:0]   _zz_addra_48;
  wire       [12:0]   _zz_addra_49;
  wire       [12:0]   _zz_addra_50;
  wire       [12:0]   _zz_addra_51;
  wire       [12:0]   _zz_addra_52;
  wire       [12:0]   _zz_addra_53;
  wire       [12:0]   _zz_addra_54;
  wire       [12:0]   _zz_addra_55;
  wire       [12:0]   _zz_addra_56;
  wire       [12:0]   _zz_addra_57;
  wire       [12:0]   _zz_addra_58;
  wire       [12:0]   _zz_addra_59;
  wire       [12:0]   _zz_addra_60;
  wire       [12:0]   _zz_addra_61;
  wire       [12:0]   _zz_addra_62;
  wire       [12:0]   _zz_addra_63;
  wire       [12:0]   _zz_addra_64;
  wire       [12:0]   _zz_addra_65;
  wire       [12:0]   _zz_addra_66;
  wire       [12:0]   _zz_addra_67;
  wire       [12:0]   _zz_addra_68;
  wire       [12:0]   _zz_addra_69;
  wire       [12:0]   _zz_addra_70;
  wire       [12:0]   _zz_addra_71;
  wire       [12:0]   _zz_addra_72;
  wire       [12:0]   _zz_addra_73;
  wire       [12:0]   _zz_addra_74;
  wire       [12:0]   _zz_addra_75;
  wire       [12:0]   _zz_addra_76;
  wire       [12:0]   _zz_addra_77;
  wire       [12:0]   _zz_addra_78;
  wire       [12:0]   _zz_addra_79;
  wire       [12:0]   _zz_addra_80;
  wire       [12:0]   _zz_addra_81;
  wire       [12:0]   _zz_addra_82;
  wire       [12:0]   _zz_addra_83;
  wire       [12:0]   _zz_addra_84;
  wire       [12:0]   _zz_addra_85;
  wire       [12:0]   _zz_addra_86;
  wire       [12:0]   _zz_addra_87;
  wire       [12:0]   _zz_addra_88;
  wire       [12:0]   _zz_addra_89;
  wire       [12:0]   _zz_addra_90;
  wire       [12:0]   _zz_addra_91;
  wire       [12:0]   _zz_addra_92;
  wire       [12:0]   _zz_addra_93;
  wire       [12:0]   _zz_addra_94;
  wire       [12:0]   _zz_addra_95;
  wire       [12:0]   _zz_addra_96;
  wire       [12:0]   _zz_addra_97;
  wire       [12:0]   _zz_addra_98;
  wire       [12:0]   _zz_addra_99;
  wire       [12:0]   _zz_addra_100;
  wire       [12:0]   _zz_addra_101;
  wire       [12:0]   _zz_addra_102;
  wire       [12:0]   _zz_addra_103;
  wire       [12:0]   _zz_addra_104;
  wire       [12:0]   _zz_addra_105;
  wire       [12:0]   _zz_addra_106;
  wire       [12:0]   _zz_addra_107;
  wire       [12:0]   _zz_addra_108;
  wire       [12:0]   _zz_addra_109;
  wire       [12:0]   _zz_addra_110;
  wire       [12:0]   _zz_addra_111;
  wire       [12:0]   _zz_addra_112;
  wire       [12:0]   _zz_addra_113;
  wire       [12:0]   _zz_addra_114;
  wire       [12:0]   _zz_addra_115;
  wire       [12:0]   _zz_addra_116;
  wire       [12:0]   _zz_addra_117;
  wire       [12:0]   _zz_addra_118;
  wire       [12:0]   _zz_addra_119;
  wire       [12:0]   _zz_addra_120;
  wire       [12:0]   _zz_addra_121;
  wire       [12:0]   _zz_addra_122;
  wire       [12:0]   _zz_addra_123;
  wire       [12:0]   _zz_addra_124;
  wire       [12:0]   _zz_addra_125;
  wire       [12:0]   _zz_addra_126;
  wire       [12:0]   _zz_addra_127;
  wire       [12:0]   _zz_addra_128;
  wire       [12:0]   _zz_addra_129;
  wire       [12:0]   _zz_addra_130;
  wire       [12:0]   _zz_addra_131;
  wire       [12:0]   _zz_addra_132;
  wire       [12:0]   _zz_addra_133;
  wire       [12:0]   _zz_addra_134;
  wire       [12:0]   _zz_addra_135;
  wire       [12:0]   _zz_addra_136;
  wire       [12:0]   _zz_addra_137;
  wire       [12:0]   _zz_addra_138;
  wire       [12:0]   _zz_addra_139;
  wire       [12:0]   _zz_addra_140;
  wire       [12:0]   _zz_addra_141;
  wire       [12:0]   _zz_addra_142;
  wire       [12:0]   _zz_addra_143;
  wire       [7:0]    _zz_when_WaCounter_l12_7;
  wire       [7:0]    _zz_when_WaCounter_l12_8;
  wire       [7:0]    _zz_when_WaCounter_l12_9;
  wire                fsm_initEnd;
  reg                 fsm_copyWeightEnd;
  wire                fsm_copyBiasEnd;
  wire                fsm_copyScaleEnd;
  wire                fsm_copyShiftEnd;
  reg        [5:0]    fsm_currentState;
  reg        [5:0]    fsm_nextState;
  wire                when_WaCounter_l17;
  reg        [2:0]    init_count;
  reg                 init_valid;
  wire                when_WaCounter_l12;
  reg        [7:0]    channelInTimes;
  reg        [11:0]   channelOutTimes;
  reg        [3:0]    copyTimes;
  wire                sData_fire;
  wire                when_WaCounter_l17_1;
  reg        [12:0]   copyWeightCnt_count;
  reg                 copyWeightCnt_valid;
  wire                when_WaCounter_l12_1;
  reg        [3:0]    copyWeightTimes_count;
  reg                 copyWeightTimes_valid;
  wire                when_WaCounter_l12_2;
  wire                sData_fire_1;
  wire                when_WaCounter_l17_2;
  reg        [7:0]    channelInCnt_count;
  reg                 channelInCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                sData_fire_2;
  wire                when_WaCounter_l17_3;
  reg        [3:0]    computeChannelOut_count;
  reg                 computeChannelOut_valid;
  wire                when_WaCounter_l12_4;
  reg        [3:0]    times_count;
  reg                 times_valid;
  wire                when_WaCounter_l12_5;
  reg        [11:0]   channelOutCnt_count;
  reg                 channelOutCnt_valid;
  wire                when_WaCounter_l12_6;
  wire                when_Weight_l250;
  wire                when_Weight_l256;
  wire                when_Weight_l260;
  wire                when_Weight_l262;
  wire                when_Weight_l268;
  reg                 weav_0_0;
  reg                 weav_0_1;
  reg                 weav_0_2;
  reg                 weav_0_3;
  reg                 weav_0_4;
  reg                 weav_0_5;
  reg                 weav_0_6;
  reg                 weav_0_7;
  reg                 weav_0_8;
  reg                 weav_0_9;
  reg                 weav_0_10;
  reg                 weav_0_11;
  reg                 weav_0_12;
  reg                 weav_0_13;
  reg                 weav_0_14;
  reg                 weav_0_15;
  reg                 weav_1_0;
  reg                 weav_1_1;
  reg                 weav_1_2;
  reg                 weav_1_3;
  reg                 weav_1_4;
  reg                 weav_1_5;
  reg                 weav_1_6;
  reg                 weav_1_7;
  reg                 weav_1_8;
  reg                 weav_1_9;
  reg                 weav_1_10;
  reg                 weav_1_11;
  reg                 weav_1_12;
  reg                 weav_1_13;
  reg                 weav_1_14;
  reg                 weav_1_15;
  reg                 weav_2_0;
  reg                 weav_2_1;
  reg                 weav_2_2;
  reg                 weav_2_3;
  reg                 weav_2_4;
  reg                 weav_2_5;
  reg                 weav_2_6;
  reg                 weav_2_7;
  reg                 weav_2_8;
  reg                 weav_2_9;
  reg                 weav_2_10;
  reg                 weav_2_11;
  reg                 weav_2_12;
  reg                 weav_2_13;
  reg                 weav_2_14;
  reg                 weav_2_15;
  reg                 weav_3_0;
  reg                 weav_3_1;
  reg                 weav_3_2;
  reg                 weav_3_3;
  reg                 weav_3_4;
  reg                 weav_3_5;
  reg                 weav_3_6;
  reg                 weav_3_7;
  reg                 weav_3_8;
  reg                 weav_3_9;
  reg                 weav_3_10;
  reg                 weav_3_11;
  reg                 weav_3_12;
  reg                 weav_3_13;
  reg                 weav_3_14;
  reg                 weav_3_15;
  reg                 weav_4_0;
  reg                 weav_4_1;
  reg                 weav_4_2;
  reg                 weav_4_3;
  reg                 weav_4_4;
  reg                 weav_4_5;
  reg                 weav_4_6;
  reg                 weav_4_7;
  reg                 weav_4_8;
  reg                 weav_4_9;
  reg                 weav_4_10;
  reg                 weav_4_11;
  reg                 weav_4_12;
  reg                 weav_4_13;
  reg                 weav_4_14;
  reg                 weav_4_15;
  reg                 weav_5_0;
  reg                 weav_5_1;
  reg                 weav_5_2;
  reg                 weav_5_3;
  reg                 weav_5_4;
  reg                 weav_5_5;
  reg                 weav_5_6;
  reg                 weav_5_7;
  reg                 weav_5_8;
  reg                 weav_5_9;
  reg                 weav_5_10;
  reg                 weav_5_11;
  reg                 weav_5_12;
  reg                 weav_5_13;
  reg                 weav_5_14;
  reg                 weav_5_15;
  reg                 weav_6_0;
  reg                 weav_6_1;
  reg                 weav_6_2;
  reg                 weav_6_3;
  reg                 weav_6_4;
  reg                 weav_6_5;
  reg                 weav_6_6;
  reg                 weav_6_7;
  reg                 weav_6_8;
  reg                 weav_6_9;
  reg                 weav_6_10;
  reg                 weav_6_11;
  reg                 weav_6_12;
  reg                 weav_6_13;
  reg                 weav_6_14;
  reg                 weav_6_15;
  reg                 weav_7_0;
  reg                 weav_7_1;
  reg                 weav_7_2;
  reg                 weav_7_3;
  reg                 weav_7_4;
  reg                 weav_7_5;
  reg                 weav_7_6;
  reg                 weav_7_7;
  reg                 weav_7_8;
  reg                 weav_7_9;
  reg                 weav_7_10;
  reg                 weav_7_11;
  reg                 weav_7_12;
  reg                 weav_7_13;
  reg                 weav_7_14;
  reg                 weav_7_15;
  reg                 weav_8_0;
  reg                 weav_8_1;
  reg                 weav_8_2;
  reg                 weav_8_3;
  reg                 weav_8_4;
  reg                 weav_8_5;
  reg                 weav_8_6;
  reg                 weav_8_7;
  reg                 weav_8_8;
  reg                 weav_8_9;
  reg                 weav_8_10;
  reg                 weav_8_11;
  reg                 weav_8_12;
  reg                 weav_8_13;
  reg                 weav_8_14;
  reg                 weav_8_15;
  wire                sData_fire_3;
  wire                when_Weight_l274;
  wire                when_Weight_l279;
  wire                when_Weight_l279_1;
  wire                when_Weight_l279_2;
  wire                when_Weight_l279_3;
  wire                when_Weight_l279_4;
  wire                when_Weight_l279_5;
  wire                when_Weight_l279_6;
  wire                when_Weight_l279_7;
  wire                when_Weight_l279_8;
  wire                when_Weight_l279_9;
  wire                when_Weight_l279_10;
  wire                when_Weight_l279_11;
  wire                when_Weight_l279_12;
  wire                when_Weight_l279_13;
  wire                when_Weight_l279_14;
  wire                when_Weight_l279_15;
  wire                when_Weight_l279_16;
  wire                when_Weight_l279_17;
  wire                when_Weight_l279_18;
  wire                when_Weight_l279_19;
  wire                when_Weight_l279_20;
  wire                when_Weight_l279_21;
  wire                when_Weight_l279_22;
  wire                when_Weight_l279_23;
  wire                when_Weight_l279_24;
  wire                when_Weight_l279_25;
  wire                when_Weight_l279_26;
  wire                when_Weight_l279_27;
  wire                when_Weight_l279_28;
  wire                when_Weight_l279_29;
  wire                when_Weight_l279_30;
  wire                when_Weight_l279_31;
  wire                when_Weight_l279_32;
  wire                when_Weight_l279_33;
  wire                when_Weight_l279_34;
  wire                when_Weight_l279_35;
  wire                when_Weight_l279_36;
  wire                when_Weight_l279_37;
  wire                when_Weight_l279_38;
  wire                when_Weight_l279_39;
  wire                when_Weight_l279_40;
  wire                when_Weight_l279_41;
  wire                when_Weight_l279_42;
  wire                when_Weight_l279_43;
  wire                when_Weight_l279_44;
  wire                when_Weight_l279_45;
  wire                when_Weight_l279_46;
  wire                when_Weight_l279_47;
  wire                when_Weight_l279_48;
  wire                when_Weight_l279_49;
  wire                when_Weight_l279_50;
  wire                when_Weight_l279_51;
  wire                when_Weight_l279_52;
  wire                when_Weight_l279_53;
  wire                when_Weight_l279_54;
  wire                when_Weight_l279_55;
  wire                when_Weight_l279_56;
  wire                when_Weight_l279_57;
  wire                when_Weight_l279_58;
  wire                when_Weight_l279_59;
  wire                when_Weight_l279_60;
  wire                when_Weight_l279_61;
  wire                when_Weight_l279_62;
  wire                when_Weight_l279_63;
  wire                when_Weight_l279_64;
  wire                when_Weight_l279_65;
  wire                when_Weight_l279_66;
  wire                when_Weight_l279_67;
  wire                when_Weight_l279_68;
  wire                when_Weight_l279_69;
  wire                when_Weight_l279_70;
  wire                when_Weight_l279_71;
  wire                when_Weight_l279_72;
  wire                when_Weight_l279_73;
  wire                when_Weight_l279_74;
  wire                when_Weight_l279_75;
  wire                when_Weight_l279_76;
  wire                when_Weight_l279_77;
  wire                when_Weight_l279_78;
  wire                when_Weight_l279_79;
  wire                when_Weight_l279_80;
  wire                when_Weight_l279_81;
  wire                when_Weight_l279_82;
  wire                when_Weight_l279_83;
  wire                when_Weight_l279_84;
  wire                when_Weight_l279_85;
  wire                when_Weight_l279_86;
  wire                when_Weight_l279_87;
  wire                when_Weight_l279_88;
  wire                when_Weight_l279_89;
  wire                when_Weight_l279_90;
  wire                when_Weight_l279_91;
  wire                when_Weight_l279_92;
  wire                when_Weight_l279_93;
  wire                when_Weight_l279_94;
  wire                when_Weight_l279_95;
  wire                when_Weight_l279_96;
  wire                when_Weight_l279_97;
  wire                when_Weight_l279_98;
  wire                when_Weight_l279_99;
  wire                when_Weight_l279_100;
  wire                when_Weight_l279_101;
  wire                when_Weight_l279_102;
  wire                when_Weight_l279_103;
  wire                when_Weight_l279_104;
  wire                when_Weight_l279_105;
  wire                when_Weight_l279_106;
  wire                when_Weight_l279_107;
  wire                when_Weight_l279_108;
  wire                when_Weight_l279_109;
  wire                when_Weight_l279_110;
  wire                when_Weight_l279_111;
  wire                when_Weight_l279_112;
  wire                when_Weight_l279_113;
  wire                when_Weight_l279_114;
  wire                when_Weight_l279_115;
  wire                when_Weight_l279_116;
  wire                when_Weight_l279_117;
  wire                when_Weight_l279_118;
  wire                when_Weight_l279_119;
  wire                when_Weight_l279_120;
  wire                when_Weight_l279_121;
  wire                when_Weight_l279_122;
  wire                when_Weight_l279_123;
  wire                when_Weight_l279_124;
  wire                when_Weight_l279_125;
  wire                when_Weight_l279_126;
  wire                when_Weight_l279_127;
  wire                when_Weight_l279_128;
  wire                when_Weight_l279_129;
  wire                when_Weight_l279_130;
  wire                when_Weight_l279_131;
  wire                when_Weight_l279_132;
  wire                when_Weight_l279_133;
  wire                when_Weight_l279_134;
  wire                when_Weight_l279_135;
  wire                when_Weight_l279_136;
  wire                when_Weight_l279_137;
  wire                when_Weight_l279_138;
  wire                when_Weight_l279_139;
  wire                when_Weight_l279_140;
  wire                when_Weight_l279_141;
  wire                when_Weight_l279_142;
  wire                when_Weight_l279_143;
  wire                when_Weight_l296;
  wire                when_Weight_l296_1;
  wire                when_Weight_l296_2;
  wire                when_Weight_l296_3;
  wire                when_Weight_l296_4;
  wire                when_Weight_l296_5;
  wire                when_Weight_l296_6;
  wire                when_Weight_l296_7;
  wire                when_Weight_l296_8;
  wire                when_Weight_l296_9;
  wire                when_Weight_l296_10;
  wire                when_Weight_l296_11;
  wire                when_Weight_l296_12;
  wire                when_Weight_l296_13;
  wire                when_Weight_l296_14;
  wire                when_Weight_l296_15;
  wire                when_Weight_l306;
  wire                when_Weight_l306_1;
  wire                when_Weight_l306_2;
  wire                when_Weight_l306_3;
  wire                when_Weight_l306_4;
  wire                when_Weight_l306_5;
  wire                when_Weight_l306_6;
  wire                when_Weight_l306_7;
  wire                when_Weight_l306_8;
  wire                when_Weight_l306_9;
  wire                when_Weight_l306_10;
  wire                when_Weight_l306_11;
  wire                when_Weight_l306_12;
  wire                when_Weight_l306_13;
  wire                when_Weight_l306_14;
  wire                when_Weight_l306_15;
  wire                when_Weight_l306_16;
  wire                when_Weight_l306_17;
  wire                when_Weight_l306_18;
  wire                when_Weight_l306_19;
  wire                when_Weight_l306_20;
  wire                when_Weight_l306_21;
  wire                when_Weight_l306_22;
  wire                when_Weight_l306_23;
  wire                when_Weight_l306_24;
  wire                when_Weight_l306_25;
  wire                when_Weight_l306_26;
  wire                when_Weight_l306_27;
  wire                when_Weight_l306_28;
  wire                when_Weight_l306_29;
  wire                when_Weight_l306_30;
  wire                when_Weight_l306_31;
  wire                when_Weight_l306_32;
  wire                when_Weight_l306_33;
  wire                when_Weight_l306_34;
  wire                when_Weight_l306_35;
  wire                when_Weight_l306_36;
  wire                when_Weight_l306_37;
  wire                when_Weight_l306_38;
  wire                when_Weight_l306_39;
  wire                when_Weight_l306_40;
  wire                when_Weight_l306_41;
  wire                when_Weight_l306_42;
  wire                when_Weight_l306_43;
  wire                when_Weight_l306_44;
  wire                when_Weight_l306_45;
  wire                when_Weight_l306_46;
  wire                when_Weight_l306_47;
  wire                when_Weight_l306_48;
  wire                when_Weight_l306_49;
  wire                when_Weight_l306_50;
  wire                when_Weight_l306_51;
  wire                when_Weight_l306_52;
  wire                when_Weight_l306_53;
  wire                when_Weight_l306_54;
  wire                when_Weight_l306_55;
  wire                when_Weight_l306_56;
  wire                when_Weight_l306_57;
  wire                when_Weight_l306_58;
  wire                when_Weight_l306_59;
  wire                when_Weight_l306_60;
  wire                when_Weight_l306_61;
  wire                when_Weight_l306_62;
  wire                when_Weight_l306_63;
  wire                when_Weight_l306_64;
  wire                when_Weight_l306_65;
  wire                when_Weight_l306_66;
  wire                when_Weight_l306_67;
  wire                when_Weight_l306_68;
  wire                when_Weight_l306_69;
  wire                when_Weight_l306_70;
  wire                when_Weight_l306_71;
  wire                when_Weight_l306_72;
  wire                when_Weight_l306_73;
  wire                when_Weight_l306_74;
  wire                when_Weight_l306_75;
  wire                when_Weight_l306_76;
  wire                when_Weight_l306_77;
  wire                when_Weight_l306_78;
  wire                when_Weight_l306_79;
  wire                when_Weight_l306_80;
  wire                when_Weight_l306_81;
  wire                when_Weight_l306_82;
  wire                when_Weight_l306_83;
  wire                when_Weight_l306_84;
  wire                when_Weight_l306_85;
  wire                when_Weight_l306_86;
  wire                when_Weight_l306_87;
  wire                when_Weight_l306_88;
  wire                when_Weight_l306_89;
  wire                when_Weight_l306_90;
  wire                when_Weight_l306_91;
  wire                when_Weight_l306_92;
  wire                when_Weight_l306_93;
  wire                when_Weight_l306_94;
  wire                when_Weight_l306_95;
  wire                when_Weight_l306_96;
  wire                when_Weight_l306_97;
  wire                when_Weight_l306_98;
  wire                when_Weight_l306_99;
  wire                when_Weight_l306_100;
  wire                when_Weight_l306_101;
  wire                when_Weight_l306_102;
  wire                when_Weight_l306_103;
  wire                when_Weight_l306_104;
  wire                when_Weight_l306_105;
  wire                when_Weight_l306_106;
  wire                when_Weight_l306_107;
  wire                when_Weight_l306_108;
  wire                when_Weight_l306_109;
  wire                when_Weight_l306_110;
  wire                when_Weight_l306_111;
  wire                when_Weight_l306_112;
  wire                when_Weight_l306_113;
  wire                when_Weight_l306_114;
  wire                when_Weight_l306_115;
  wire                when_Weight_l306_116;
  wire                when_Weight_l306_117;
  wire                when_Weight_l306_118;
  wire                when_Weight_l306_119;
  wire                when_Weight_l306_120;
  wire                when_Weight_l306_121;
  wire                when_Weight_l306_122;
  wire                when_Weight_l306_123;
  wire                when_Weight_l306_124;
  wire                when_Weight_l306_125;
  wire                when_Weight_l306_126;
  wire                when_Weight_l306_127;
  reg        [12:0]   addr_0_0;
  reg        [12:0]   addr_0_1;
  reg        [12:0]   addr_0_2;
  reg        [12:0]   addr_0_3;
  reg        [12:0]   addr_0_4;
  reg        [12:0]   addr_0_5;
  reg        [12:0]   addr_0_6;
  reg        [12:0]   addr_0_7;
  reg        [12:0]   addr_0_8;
  reg        [12:0]   addr_0_9;
  reg        [12:0]   addr_0_10;
  reg        [12:0]   addr_0_11;
  reg        [12:0]   addr_0_12;
  reg        [12:0]   addr_0_13;
  reg        [12:0]   addr_0_14;
  reg        [12:0]   addr_0_15;
  reg        [12:0]   addr_1_0;
  reg        [12:0]   addr_1_1;
  reg        [12:0]   addr_1_2;
  reg        [12:0]   addr_1_3;
  reg        [12:0]   addr_1_4;
  reg        [12:0]   addr_1_5;
  reg        [12:0]   addr_1_6;
  reg        [12:0]   addr_1_7;
  reg        [12:0]   addr_1_8;
  reg        [12:0]   addr_1_9;
  reg        [12:0]   addr_1_10;
  reg        [12:0]   addr_1_11;
  reg        [12:0]   addr_1_12;
  reg        [12:0]   addr_1_13;
  reg        [12:0]   addr_1_14;
  reg        [12:0]   addr_1_15;
  reg        [12:0]   addr_2_0;
  reg        [12:0]   addr_2_1;
  reg        [12:0]   addr_2_2;
  reg        [12:0]   addr_2_3;
  reg        [12:0]   addr_2_4;
  reg        [12:0]   addr_2_5;
  reg        [12:0]   addr_2_6;
  reg        [12:0]   addr_2_7;
  reg        [12:0]   addr_2_8;
  reg        [12:0]   addr_2_9;
  reg        [12:0]   addr_2_10;
  reg        [12:0]   addr_2_11;
  reg        [12:0]   addr_2_12;
  reg        [12:0]   addr_2_13;
  reg        [12:0]   addr_2_14;
  reg        [12:0]   addr_2_15;
  reg        [12:0]   addr_3_0;
  reg        [12:0]   addr_3_1;
  reg        [12:0]   addr_3_2;
  reg        [12:0]   addr_3_3;
  reg        [12:0]   addr_3_4;
  reg        [12:0]   addr_3_5;
  reg        [12:0]   addr_3_6;
  reg        [12:0]   addr_3_7;
  reg        [12:0]   addr_3_8;
  reg        [12:0]   addr_3_9;
  reg        [12:0]   addr_3_10;
  reg        [12:0]   addr_3_11;
  reg        [12:0]   addr_3_12;
  reg        [12:0]   addr_3_13;
  reg        [12:0]   addr_3_14;
  reg        [12:0]   addr_3_15;
  reg        [12:0]   addr_4_0;
  reg        [12:0]   addr_4_1;
  reg        [12:0]   addr_4_2;
  reg        [12:0]   addr_4_3;
  reg        [12:0]   addr_4_4;
  reg        [12:0]   addr_4_5;
  reg        [12:0]   addr_4_6;
  reg        [12:0]   addr_4_7;
  reg        [12:0]   addr_4_8;
  reg        [12:0]   addr_4_9;
  reg        [12:0]   addr_4_10;
  reg        [12:0]   addr_4_11;
  reg        [12:0]   addr_4_12;
  reg        [12:0]   addr_4_13;
  reg        [12:0]   addr_4_14;
  reg        [12:0]   addr_4_15;
  reg        [12:0]   addr_5_0;
  reg        [12:0]   addr_5_1;
  reg        [12:0]   addr_5_2;
  reg        [12:0]   addr_5_3;
  reg        [12:0]   addr_5_4;
  reg        [12:0]   addr_5_5;
  reg        [12:0]   addr_5_6;
  reg        [12:0]   addr_5_7;
  reg        [12:0]   addr_5_8;
  reg        [12:0]   addr_5_9;
  reg        [12:0]   addr_5_10;
  reg        [12:0]   addr_5_11;
  reg        [12:0]   addr_5_12;
  reg        [12:0]   addr_5_13;
  reg        [12:0]   addr_5_14;
  reg        [12:0]   addr_5_15;
  reg        [12:0]   addr_6_0;
  reg        [12:0]   addr_6_1;
  reg        [12:0]   addr_6_2;
  reg        [12:0]   addr_6_3;
  reg        [12:0]   addr_6_4;
  reg        [12:0]   addr_6_5;
  reg        [12:0]   addr_6_6;
  reg        [12:0]   addr_6_7;
  reg        [12:0]   addr_6_8;
  reg        [12:0]   addr_6_9;
  reg        [12:0]   addr_6_10;
  reg        [12:0]   addr_6_11;
  reg        [12:0]   addr_6_12;
  reg        [12:0]   addr_6_13;
  reg        [12:0]   addr_6_14;
  reg        [12:0]   addr_6_15;
  reg        [12:0]   addr_7_0;
  reg        [12:0]   addr_7_1;
  reg        [12:0]   addr_7_2;
  reg        [12:0]   addr_7_3;
  reg        [12:0]   addr_7_4;
  reg        [12:0]   addr_7_5;
  reg        [12:0]   addr_7_6;
  reg        [12:0]   addr_7_7;
  reg        [12:0]   addr_7_8;
  reg        [12:0]   addr_7_9;
  reg        [12:0]   addr_7_10;
  reg        [12:0]   addr_7_11;
  reg        [12:0]   addr_7_12;
  reg        [12:0]   addr_7_13;
  reg        [12:0]   addr_7_14;
  reg        [12:0]   addr_7_15;
  reg        [12:0]   addr_8_0;
  reg        [12:0]   addr_8_1;
  reg        [12:0]   addr_8_2;
  reg        [12:0]   addr_8_3;
  reg        [12:0]   addr_8_4;
  reg        [12:0]   addr_8_5;
  reg        [12:0]   addr_8_6;
  reg        [12:0]   addr_8_7;
  reg        [12:0]   addr_8_8;
  reg        [12:0]   addr_8_9;
  reg        [12:0]   addr_8_10;
  reg        [12:0]   addr_8_11;
  reg        [12:0]   addr_8_12;
  reg        [12:0]   addr_8_13;
  reg        [12:0]   addr_8_14;
  reg        [12:0]   addr_8_15;
  wire                when_Weight_l326;
  wire                when_Weight_l326_1;
  wire                when_Weight_l326_2;
  wire                when_Weight_l326_3;
  wire                when_Weight_l326_4;
  wire                when_Weight_l326_5;
  wire                when_Weight_l326_6;
  wire                when_Weight_l326_7;
  wire                when_Weight_l326_8;
  wire                when_Weight_l326_9;
  wire                when_Weight_l326_10;
  wire                when_Weight_l326_11;
  wire                when_Weight_l326_12;
  wire                when_Weight_l326_13;
  wire                when_Weight_l326_14;
  wire                when_Weight_l326_15;
  wire                when_Weight_l326_16;
  wire                when_Weight_l326_17;
  wire                when_Weight_l326_18;
  wire                when_Weight_l326_19;
  wire                when_Weight_l326_20;
  wire                when_Weight_l326_21;
  wire                when_Weight_l326_22;
  wire                when_Weight_l326_23;
  wire                when_Weight_l326_24;
  wire                when_Weight_l326_25;
  wire                when_Weight_l326_26;
  wire                when_Weight_l326_27;
  wire                when_Weight_l326_28;
  wire                when_Weight_l326_29;
  wire                when_Weight_l326_30;
  wire                when_Weight_l326_31;
  wire                when_Weight_l326_32;
  wire                when_Weight_l326_33;
  wire                when_Weight_l326_34;
  wire                when_Weight_l326_35;
  wire                when_Weight_l326_36;
  wire                when_Weight_l326_37;
  wire                when_Weight_l326_38;
  wire                when_Weight_l326_39;
  wire                when_Weight_l326_40;
  wire                when_Weight_l326_41;
  wire                when_Weight_l326_42;
  wire                when_Weight_l326_43;
  wire                when_Weight_l326_44;
  wire                when_Weight_l326_45;
  wire                when_Weight_l326_46;
  wire                when_Weight_l326_47;
  wire                when_Weight_l326_48;
  wire                when_Weight_l326_49;
  wire                when_Weight_l326_50;
  wire                when_Weight_l326_51;
  wire                when_Weight_l326_52;
  wire                when_Weight_l326_53;
  wire                when_Weight_l326_54;
  wire                when_Weight_l326_55;
  wire                when_Weight_l326_56;
  wire                when_Weight_l326_57;
  wire                when_Weight_l326_58;
  wire                when_Weight_l326_59;
  wire                when_Weight_l326_60;
  wire                when_Weight_l326_61;
  wire                when_Weight_l326_62;
  wire                when_Weight_l326_63;
  wire                when_Weight_l326_64;
  wire                when_Weight_l326_65;
  wire                when_Weight_l326_66;
  wire                when_Weight_l326_67;
  wire                when_Weight_l326_68;
  wire                when_Weight_l326_69;
  wire                when_Weight_l326_70;
  wire                when_Weight_l326_71;
  wire                when_Weight_l326_72;
  wire                when_Weight_l326_73;
  wire                when_Weight_l326_74;
  wire                when_Weight_l326_75;
  wire                when_Weight_l326_76;
  wire                when_Weight_l326_77;
  wire                when_Weight_l326_78;
  wire                when_Weight_l326_79;
  wire                when_Weight_l326_80;
  wire                when_Weight_l326_81;
  wire                when_Weight_l326_82;
  wire                when_Weight_l326_83;
  wire                when_Weight_l326_84;
  wire                when_Weight_l326_85;
  wire                when_Weight_l326_86;
  wire                when_Weight_l326_87;
  wire                when_Weight_l326_88;
  wire                when_Weight_l326_89;
  wire                when_Weight_l326_90;
  wire                when_Weight_l326_91;
  wire                when_Weight_l326_92;
  wire                when_Weight_l326_93;
  wire                when_Weight_l326_94;
  wire                when_Weight_l326_95;
  wire                when_Weight_l326_96;
  wire                when_Weight_l326_97;
  wire                when_Weight_l326_98;
  wire                when_Weight_l326_99;
  wire                when_Weight_l326_100;
  wire                when_Weight_l326_101;
  wire                when_Weight_l326_102;
  wire                when_Weight_l326_103;
  wire                when_Weight_l326_104;
  wire                when_Weight_l326_105;
  wire                when_Weight_l326_106;
  wire                when_Weight_l326_107;
  wire                when_Weight_l326_108;
  wire                when_Weight_l326_109;
  wire                when_Weight_l326_110;
  wire                when_Weight_l326_111;
  wire                when_Weight_l326_112;
  wire                when_Weight_l326_113;
  wire                when_Weight_l326_114;
  wire                when_Weight_l326_115;
  wire                when_Weight_l326_116;
  wire                when_Weight_l326_117;
  wire                when_Weight_l326_118;
  wire                when_Weight_l326_119;
  wire                when_Weight_l326_120;
  wire                when_Weight_l326_121;
  wire                when_Weight_l326_122;
  wire                when_Weight_l326_123;
  wire                when_Weight_l326_124;
  wire                when_Weight_l326_125;
  wire                when_Weight_l326_126;
  wire                when_Weight_l326_127;
  wire                when_Weight_l326_128;
  wire                when_Weight_l326_129;
  wire                when_Weight_l326_130;
  wire                when_Weight_l326_131;
  wire                when_Weight_l326_132;
  wire                when_Weight_l326_133;
  wire                when_Weight_l326_134;
  wire                when_Weight_l326_135;
  wire                when_Weight_l326_136;
  wire                when_Weight_l326_137;
  wire                when_Weight_l326_138;
  wire                when_Weight_l326_139;
  wire                when_Weight_l326_140;
  wire                when_Weight_l326_141;
  wire                when_Weight_l326_142;
  wire                when_Weight_l326_143;
  wire       [127:0]  weightData_0_0;
  wire       [127:0]  weightData_0_1;
  wire       [127:0]  weightData_0_2;
  wire       [127:0]  weightData_0_3;
  wire       [127:0]  weightData_0_4;
  wire       [127:0]  weightData_0_5;
  wire       [127:0]  weightData_0_6;
  wire       [127:0]  weightData_0_7;
  wire       [127:0]  weightData_0_8;
  wire       [127:0]  weightData_0_9;
  wire       [127:0]  weightData_0_10;
  wire       [127:0]  weightData_0_11;
  wire       [127:0]  weightData_0_12;
  wire       [127:0]  weightData_0_13;
  wire       [127:0]  weightData_0_14;
  wire       [127:0]  weightData_0_15;
  wire       [127:0]  weightData_1_0;
  wire       [127:0]  weightData_1_1;
  wire       [127:0]  weightData_1_2;
  wire       [127:0]  weightData_1_3;
  wire       [127:0]  weightData_1_4;
  wire       [127:0]  weightData_1_5;
  wire       [127:0]  weightData_1_6;
  wire       [127:0]  weightData_1_7;
  wire       [127:0]  weightData_1_8;
  wire       [127:0]  weightData_1_9;
  wire       [127:0]  weightData_1_10;
  wire       [127:0]  weightData_1_11;
  wire       [127:0]  weightData_1_12;
  wire       [127:0]  weightData_1_13;
  wire       [127:0]  weightData_1_14;
  wire       [127:0]  weightData_1_15;
  wire       [127:0]  weightData_2_0;
  wire       [127:0]  weightData_2_1;
  wire       [127:0]  weightData_2_2;
  wire       [127:0]  weightData_2_3;
  wire       [127:0]  weightData_2_4;
  wire       [127:0]  weightData_2_5;
  wire       [127:0]  weightData_2_6;
  wire       [127:0]  weightData_2_7;
  wire       [127:0]  weightData_2_8;
  wire       [127:0]  weightData_2_9;
  wire       [127:0]  weightData_2_10;
  wire       [127:0]  weightData_2_11;
  wire       [127:0]  weightData_2_12;
  wire       [127:0]  weightData_2_13;
  wire       [127:0]  weightData_2_14;
  wire       [127:0]  weightData_2_15;
  wire       [127:0]  weightData_3_0;
  wire       [127:0]  weightData_3_1;
  wire       [127:0]  weightData_3_2;
  wire       [127:0]  weightData_3_3;
  wire       [127:0]  weightData_3_4;
  wire       [127:0]  weightData_3_5;
  wire       [127:0]  weightData_3_6;
  wire       [127:0]  weightData_3_7;
  wire       [127:0]  weightData_3_8;
  wire       [127:0]  weightData_3_9;
  wire       [127:0]  weightData_3_10;
  wire       [127:0]  weightData_3_11;
  wire       [127:0]  weightData_3_12;
  wire       [127:0]  weightData_3_13;
  wire       [127:0]  weightData_3_14;
  wire       [127:0]  weightData_3_15;
  wire       [127:0]  weightData_4_0;
  wire       [127:0]  weightData_4_1;
  wire       [127:0]  weightData_4_2;
  wire       [127:0]  weightData_4_3;
  wire       [127:0]  weightData_4_4;
  wire       [127:0]  weightData_4_5;
  wire       [127:0]  weightData_4_6;
  wire       [127:0]  weightData_4_7;
  wire       [127:0]  weightData_4_8;
  wire       [127:0]  weightData_4_9;
  wire       [127:0]  weightData_4_10;
  wire       [127:0]  weightData_4_11;
  wire       [127:0]  weightData_4_12;
  wire       [127:0]  weightData_4_13;
  wire       [127:0]  weightData_4_14;
  wire       [127:0]  weightData_4_15;
  wire       [127:0]  weightData_5_0;
  wire       [127:0]  weightData_5_1;
  wire       [127:0]  weightData_5_2;
  wire       [127:0]  weightData_5_3;
  wire       [127:0]  weightData_5_4;
  wire       [127:0]  weightData_5_5;
  wire       [127:0]  weightData_5_6;
  wire       [127:0]  weightData_5_7;
  wire       [127:0]  weightData_5_8;
  wire       [127:0]  weightData_5_9;
  wire       [127:0]  weightData_5_10;
  wire       [127:0]  weightData_5_11;
  wire       [127:0]  weightData_5_12;
  wire       [127:0]  weightData_5_13;
  wire       [127:0]  weightData_5_14;
  wire       [127:0]  weightData_5_15;
  wire       [127:0]  weightData_6_0;
  wire       [127:0]  weightData_6_1;
  wire       [127:0]  weightData_6_2;
  wire       [127:0]  weightData_6_3;
  wire       [127:0]  weightData_6_4;
  wire       [127:0]  weightData_6_5;
  wire       [127:0]  weightData_6_6;
  wire       [127:0]  weightData_6_7;
  wire       [127:0]  weightData_6_8;
  wire       [127:0]  weightData_6_9;
  wire       [127:0]  weightData_6_10;
  wire       [127:0]  weightData_6_11;
  wire       [127:0]  weightData_6_12;
  wire       [127:0]  weightData_6_13;
  wire       [127:0]  weightData_6_14;
  wire       [127:0]  weightData_6_15;
  wire       [127:0]  weightData_7_0;
  wire       [127:0]  weightData_7_1;
  wire       [127:0]  weightData_7_2;
  wire       [127:0]  weightData_7_3;
  wire       [127:0]  weightData_7_4;
  wire       [127:0]  weightData_7_5;
  wire       [127:0]  weightData_7_6;
  wire       [127:0]  weightData_7_7;
  wire       [127:0]  weightData_7_8;
  wire       [127:0]  weightData_7_9;
  wire       [127:0]  weightData_7_10;
  wire       [127:0]  weightData_7_11;
  wire       [127:0]  weightData_7_12;
  wire       [127:0]  weightData_7_13;
  wire       [127:0]  weightData_7_14;
  wire       [127:0]  weightData_7_15;
  wire       [127:0]  weightData_8_0;
  wire       [127:0]  weightData_8_1;
  wire       [127:0]  weightData_8_2;
  wire       [127:0]  weightData_8_3;
  wire       [127:0]  weightData_8_4;
  wire       [127:0]  weightData_8_5;
  wire       [127:0]  weightData_8_6;
  wire       [127:0]  weightData_8_7;
  wire       [127:0]  weightData_8_8;
  wire       [127:0]  weightData_8_9;
  wire       [127:0]  weightData_8_10;
  wire       [127:0]  weightData_8_11;
  wire       [127:0]  weightData_8_12;
  wire       [127:0]  weightData_8_13;
  wire       [127:0]  weightData_8_14;
  wire       [127:0]  weightData_8_15;
  wire                sData_fire_4;
  wire                when_WaCounter_l17_4;
  wire                sData_fire_5;
  reg        [7:0]    copyBias_copyCnt_count;
  reg                 copyBias_copyCnt_valid;
  wire                when_WaCounter_l12_7;
  wire                sData_fire_6;
  wire                when_WaCounter_l17_5;
  wire                sData_fire_7;
  reg        [7:0]    copyScale_copyCnt_count;
  reg                 copyScale_copyCnt_valid;
  wire                when_WaCounter_l12_8;
  wire                sData_fire_8;
  wire                when_WaCounter_l17_6;
  wire                sData_fire_9;
  reg        [7:0]    copyShift_copyCnt_count;
  reg                 copyShift_copyCnt_valid;
  wire                when_WaCounter_l12_9;
  wire                when_WaUtil_l29;
  `ifndef SYNTHESIS
  reg [87:0] fsm_currentState_string;
  reg [87:0] fsm_nextState_string;
  `endif


  assign _zz_when_WaCounter_l12_1 = (weightNum - 13'h0001);
  assign _zz_when_WaCounter_l12_3 = (channelInTimes - 8'h01);
  assign _zz_when_WaCounter_l12_6 = (channelOutTimes - 12'h001);
  assign _zz_when_Weight_l326 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_1 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_2 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_3 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_4 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_5 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_6 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_7 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_8 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_9 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_10 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_11 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_12 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_13 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_14 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_15 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_16 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_17 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_18 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_19 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_20 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_21 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_22 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_23 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_24 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_25 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_26 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_27 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_28 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_29 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_30 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_31 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_32 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_33 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_34 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_35 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_36 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_37 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_38 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_39 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_40 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_41 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_42 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_43 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_44 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_45 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_46 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_47 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_48 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_49 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_50 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_51 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_52 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_53 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_54 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_55 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_56 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_57 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_58 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_59 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_60 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_61 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_62 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_63 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_64 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_65 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_66 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_67 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_68 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_69 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_70 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_71 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_72 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_73 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_74 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_75 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_76 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_77 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_78 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_79 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_80 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_81 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_82 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_83 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_84 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_85 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_86 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_87 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_88 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_89 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_90 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_91 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_92 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_93 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_94 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_95 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_96 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_97 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_98 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_99 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_100 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_101 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_102 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_103 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_104 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_105 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_106 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_107 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_108 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_109 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_110 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_111 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_112 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_113 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_114 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_115 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_116 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_117 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_118 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_119 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_120 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_121 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_122 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_123 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_124 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_125 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_126 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_127 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_128 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_129 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_130 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_131 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_132 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_133 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_134 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_135 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_136 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_137 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_138 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_139 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_140 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_141 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_142 = (weightNum - 13'h0001);
  assign _zz_when_Weight_l326_143 = (weightNum - 13'h0001);
  assign _zz_addra = addr_0_0;
  assign _zz_addra_1 = addr_0_1;
  assign _zz_addra_2 = addr_0_2;
  assign _zz_addra_3 = addr_0_3;
  assign _zz_addra_4 = addr_0_4;
  assign _zz_addra_5 = addr_0_5;
  assign _zz_addra_6 = addr_0_6;
  assign _zz_addra_7 = addr_0_7;
  assign _zz_addra_8 = addr_0_8;
  assign _zz_addra_9 = addr_0_9;
  assign _zz_addra_10 = addr_0_10;
  assign _zz_addra_11 = addr_0_11;
  assign _zz_addra_12 = addr_0_12;
  assign _zz_addra_13 = addr_0_13;
  assign _zz_addra_14 = addr_0_14;
  assign _zz_addra_15 = addr_0_15;
  assign _zz_addra_16 = addr_1_0;
  assign _zz_addra_17 = addr_1_1;
  assign _zz_addra_18 = addr_1_2;
  assign _zz_addra_19 = addr_1_3;
  assign _zz_addra_20 = addr_1_4;
  assign _zz_addra_21 = addr_1_5;
  assign _zz_addra_22 = addr_1_6;
  assign _zz_addra_23 = addr_1_7;
  assign _zz_addra_24 = addr_1_8;
  assign _zz_addra_25 = addr_1_9;
  assign _zz_addra_26 = addr_1_10;
  assign _zz_addra_27 = addr_1_11;
  assign _zz_addra_28 = addr_1_12;
  assign _zz_addra_29 = addr_1_13;
  assign _zz_addra_30 = addr_1_14;
  assign _zz_addra_31 = addr_1_15;
  assign _zz_addra_32 = addr_2_0;
  assign _zz_addra_33 = addr_2_1;
  assign _zz_addra_34 = addr_2_2;
  assign _zz_addra_35 = addr_2_3;
  assign _zz_addra_36 = addr_2_4;
  assign _zz_addra_37 = addr_2_5;
  assign _zz_addra_38 = addr_2_6;
  assign _zz_addra_39 = addr_2_7;
  assign _zz_addra_40 = addr_2_8;
  assign _zz_addra_41 = addr_2_9;
  assign _zz_addra_42 = addr_2_10;
  assign _zz_addra_43 = addr_2_11;
  assign _zz_addra_44 = addr_2_12;
  assign _zz_addra_45 = addr_2_13;
  assign _zz_addra_46 = addr_2_14;
  assign _zz_addra_47 = addr_2_15;
  assign _zz_addra_48 = addr_3_0;
  assign _zz_addra_49 = addr_3_1;
  assign _zz_addra_50 = addr_3_2;
  assign _zz_addra_51 = addr_3_3;
  assign _zz_addra_52 = addr_3_4;
  assign _zz_addra_53 = addr_3_5;
  assign _zz_addra_54 = addr_3_6;
  assign _zz_addra_55 = addr_3_7;
  assign _zz_addra_56 = addr_3_8;
  assign _zz_addra_57 = addr_3_9;
  assign _zz_addra_58 = addr_3_10;
  assign _zz_addra_59 = addr_3_11;
  assign _zz_addra_60 = addr_3_12;
  assign _zz_addra_61 = addr_3_13;
  assign _zz_addra_62 = addr_3_14;
  assign _zz_addra_63 = addr_3_15;
  assign _zz_addra_64 = addr_4_0;
  assign _zz_addra_65 = addr_4_1;
  assign _zz_addra_66 = addr_4_2;
  assign _zz_addra_67 = addr_4_3;
  assign _zz_addra_68 = addr_4_4;
  assign _zz_addra_69 = addr_4_5;
  assign _zz_addra_70 = addr_4_6;
  assign _zz_addra_71 = addr_4_7;
  assign _zz_addra_72 = addr_4_8;
  assign _zz_addra_73 = addr_4_9;
  assign _zz_addra_74 = addr_4_10;
  assign _zz_addra_75 = addr_4_11;
  assign _zz_addra_76 = addr_4_12;
  assign _zz_addra_77 = addr_4_13;
  assign _zz_addra_78 = addr_4_14;
  assign _zz_addra_79 = addr_4_15;
  assign _zz_addra_80 = addr_5_0;
  assign _zz_addra_81 = addr_5_1;
  assign _zz_addra_82 = addr_5_2;
  assign _zz_addra_83 = addr_5_3;
  assign _zz_addra_84 = addr_5_4;
  assign _zz_addra_85 = addr_5_5;
  assign _zz_addra_86 = addr_5_6;
  assign _zz_addra_87 = addr_5_7;
  assign _zz_addra_88 = addr_5_8;
  assign _zz_addra_89 = addr_5_9;
  assign _zz_addra_90 = addr_5_10;
  assign _zz_addra_91 = addr_5_11;
  assign _zz_addra_92 = addr_5_12;
  assign _zz_addra_93 = addr_5_13;
  assign _zz_addra_94 = addr_5_14;
  assign _zz_addra_95 = addr_5_15;
  assign _zz_addra_96 = addr_6_0;
  assign _zz_addra_97 = addr_6_1;
  assign _zz_addra_98 = addr_6_2;
  assign _zz_addra_99 = addr_6_3;
  assign _zz_addra_100 = addr_6_4;
  assign _zz_addra_101 = addr_6_5;
  assign _zz_addra_102 = addr_6_6;
  assign _zz_addra_103 = addr_6_7;
  assign _zz_addra_104 = addr_6_8;
  assign _zz_addra_105 = addr_6_9;
  assign _zz_addra_106 = addr_6_10;
  assign _zz_addra_107 = addr_6_11;
  assign _zz_addra_108 = addr_6_12;
  assign _zz_addra_109 = addr_6_13;
  assign _zz_addra_110 = addr_6_14;
  assign _zz_addra_111 = addr_6_15;
  assign _zz_addra_112 = addr_7_0;
  assign _zz_addra_113 = addr_7_1;
  assign _zz_addra_114 = addr_7_2;
  assign _zz_addra_115 = addr_7_3;
  assign _zz_addra_116 = addr_7_4;
  assign _zz_addra_117 = addr_7_5;
  assign _zz_addra_118 = addr_7_6;
  assign _zz_addra_119 = addr_7_7;
  assign _zz_addra_120 = addr_7_8;
  assign _zz_addra_121 = addr_7_9;
  assign _zz_addra_122 = addr_7_10;
  assign _zz_addra_123 = addr_7_11;
  assign _zz_addra_124 = addr_7_12;
  assign _zz_addra_125 = addr_7_13;
  assign _zz_addra_126 = addr_7_14;
  assign _zz_addra_127 = addr_7_15;
  assign _zz_addra_128 = addr_8_0;
  assign _zz_addra_129 = addr_8_1;
  assign _zz_addra_130 = addr_8_2;
  assign _zz_addra_131 = addr_8_3;
  assign _zz_addra_132 = addr_8_4;
  assign _zz_addra_133 = addr_8_5;
  assign _zz_addra_134 = addr_8_6;
  assign _zz_addra_135 = addr_8_7;
  assign _zz_addra_136 = addr_8_8;
  assign _zz_addra_137 = addr_8_9;
  assign _zz_addra_138 = addr_8_10;
  assign _zz_addra_139 = addr_8_11;
  assign _zz_addra_140 = addr_8_12;
  assign _zz_addra_141 = addr_8_13;
  assign _zz_addra_142 = addr_8_14;
  assign _zz_addra_143 = addr_8_15;
  assign _zz_when_WaCounter_l12_7 = (quanNum - 8'h01);
  assign _zz_when_WaCounter_l12_8 = (quanNum - 8'h01);
  assign _zz_when_WaCounter_l12_9 = (quanNum - 8'h01);
  assign _zz_weightRead_0_data = {{{{{{{_zz_weightRead_0_data_1,_zz_weightRead_0_data_2},weightData_0_11},weightData_0_10},weightData_0_9},weightData_0_8},weightData_0_7},weightData_0_6};
  assign _zz_weightRead_0_data_1 = {{weightData_0_15,weightData_0_14},weightData_0_13};
  assign _zz_weightRead_0_data_2 = weightData_0_12;
  assign _zz_weightRead_1_data = {{{{{{{_zz_weightRead_1_data_1,_zz_weightRead_1_data_2},weightData_1_11},weightData_1_10},weightData_1_9},weightData_1_8},weightData_1_7},weightData_1_6};
  assign _zz_weightRead_1_data_1 = {{weightData_1_15,weightData_1_14},weightData_1_13};
  assign _zz_weightRead_1_data_2 = weightData_1_12;
  assign _zz_weightRead_2_data = {{{{{{{_zz_weightRead_2_data_1,_zz_weightRead_2_data_2},weightData_2_11},weightData_2_10},weightData_2_9},weightData_2_8},weightData_2_7},weightData_2_6};
  assign _zz_weightRead_2_data_1 = {{weightData_2_15,weightData_2_14},weightData_2_13};
  assign _zz_weightRead_2_data_2 = weightData_2_12;
  assign _zz_weightRead_3_data = {{{{{{{_zz_weightRead_3_data_1,_zz_weightRead_3_data_2},weightData_3_11},weightData_3_10},weightData_3_9},weightData_3_8},weightData_3_7},weightData_3_6};
  assign _zz_weightRead_3_data_1 = {{weightData_3_15,weightData_3_14},weightData_3_13};
  assign _zz_weightRead_3_data_2 = weightData_3_12;
  assign _zz_weightRead_4_data = {{{{{{{_zz_weightRead_4_data_1,_zz_weightRead_4_data_2},weightData_4_11},weightData_4_10},weightData_4_9},weightData_4_8},weightData_4_7},weightData_4_6};
  assign _zz_weightRead_4_data_1 = {{weightData_4_15,weightData_4_14},weightData_4_13};
  assign _zz_weightRead_4_data_2 = weightData_4_12;
  assign _zz_weightRead_5_data = {{{{{{{_zz_weightRead_5_data_1,_zz_weightRead_5_data_2},weightData_5_11},weightData_5_10},weightData_5_9},weightData_5_8},weightData_5_7},weightData_5_6};
  assign _zz_weightRead_5_data_1 = {{weightData_5_15,weightData_5_14},weightData_5_13};
  assign _zz_weightRead_5_data_2 = weightData_5_12;
  assign _zz_weightRead_6_data = {{{{{{{_zz_weightRead_6_data_1,_zz_weightRead_6_data_2},weightData_6_11},weightData_6_10},weightData_6_9},weightData_6_8},weightData_6_7},weightData_6_6};
  assign _zz_weightRead_6_data_1 = {{weightData_6_15,weightData_6_14},weightData_6_13};
  assign _zz_weightRead_6_data_2 = weightData_6_12;
  assign _zz_weightRead_7_data = {{{{{{{_zz_weightRead_7_data_1,_zz_weightRead_7_data_2},weightData_7_11},weightData_7_10},weightData_7_9},weightData_7_8},weightData_7_7},weightData_7_6};
  assign _zz_weightRead_7_data_1 = {{weightData_7_15,weightData_7_14},weightData_7_13};
  assign _zz_weightRead_7_data_2 = weightData_7_12;
  assign _zz_weightRead_8_data = {{{{{{{_zz_weightRead_8_data_1,_zz_weightRead_8_data_2},weightData_8_11},weightData_8_10},weightData_8_9},weightData_8_8},weightData_8_7},weightData_8_6};
  assign _zz_weightRead_8_data_1 = {{weightData_8_15,weightData_8_14},weightData_8_13};
  assign _zz_weightRead_8_data_2 = weightData_8_12;
  sdpram weightRam_0_0 (
    .doutb (weightRam_0_0_doutb[127:0]), //o
    .addra (weightRam_0_0_addra[8:0]  ), //i
    .addrb (weightRam_0_0_addrb[8:0]  ), //i
    .dina  (weightRam_0_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_1 (
    .doutb (weightRam_0_1_doutb[127:0]), //o
    .addra (weightRam_0_1_addra[8:0]  ), //i
    .addrb (weightRam_0_1_addrb[8:0]  ), //i
    .dina  (weightRam_0_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_2 (
    .doutb (weightRam_0_2_doutb[127:0]), //o
    .addra (weightRam_0_2_addra[8:0]  ), //i
    .addrb (weightRam_0_2_addrb[8:0]  ), //i
    .dina  (weightRam_0_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_3 (
    .doutb (weightRam_0_3_doutb[127:0]), //o
    .addra (weightRam_0_3_addra[8:0]  ), //i
    .addrb (weightRam_0_3_addrb[8:0]  ), //i
    .dina  (weightRam_0_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_4 (
    .doutb (weightRam_0_4_doutb[127:0]), //o
    .addra (weightRam_0_4_addra[8:0]  ), //i
    .addrb (weightRam_0_4_addrb[8:0]  ), //i
    .dina  (weightRam_0_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_5 (
    .doutb (weightRam_0_5_doutb[127:0]), //o
    .addra (weightRam_0_5_addra[8:0]  ), //i
    .addrb (weightRam_0_5_addrb[8:0]  ), //i
    .dina  (weightRam_0_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_6 (
    .doutb (weightRam_0_6_doutb[127:0]), //o
    .addra (weightRam_0_6_addra[8:0]  ), //i
    .addrb (weightRam_0_6_addrb[8:0]  ), //i
    .dina  (weightRam_0_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_7 (
    .doutb (weightRam_0_7_doutb[127:0]), //o
    .addra (weightRam_0_7_addra[8:0]  ), //i
    .addrb (weightRam_0_7_addrb[8:0]  ), //i
    .dina  (weightRam_0_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_8 (
    .doutb (weightRam_0_8_doutb[127:0]), //o
    .addra (weightRam_0_8_addra[8:0]  ), //i
    .addrb (weightRam_0_8_addrb[8:0]  ), //i
    .dina  (weightRam_0_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_9 (
    .doutb (weightRam_0_9_doutb[127:0]), //o
    .addra (weightRam_0_9_addra[8:0]  ), //i
    .addrb (weightRam_0_9_addrb[8:0]  ), //i
    .dina  (weightRam_0_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_0_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_0_10 (
    .doutb (weightRam_0_10_doutb[127:0]), //o
    .addra (weightRam_0_10_addra[8:0]  ), //i
    .addrb (weightRam_0_10_addrb[8:0]  ), //i
    .dina  (weightRam_0_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_0_11 (
    .doutb (weightRam_0_11_doutb[127:0]), //o
    .addra (weightRam_0_11_addra[8:0]  ), //i
    .addrb (weightRam_0_11_addrb[8:0]  ), //i
    .dina  (weightRam_0_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_0_12 (
    .doutb (weightRam_0_12_doutb[127:0]), //o
    .addra (weightRam_0_12_addra[8:0]  ), //i
    .addrb (weightRam_0_12_addrb[8:0]  ), //i
    .dina  (weightRam_0_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_0_13 (
    .doutb (weightRam_0_13_doutb[127:0]), //o
    .addra (weightRam_0_13_addra[8:0]  ), //i
    .addrb (weightRam_0_13_addrb[8:0]  ), //i
    .dina  (weightRam_0_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_0_14 (
    .doutb (weightRam_0_14_doutb[127:0]), //o
    .addra (weightRam_0_14_addra[8:0]  ), //i
    .addrb (weightRam_0_14_addrb[8:0]  ), //i
    .dina  (weightRam_0_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_0_15 (
    .doutb (weightRam_0_15_doutb[127:0]), //o
    .addra (weightRam_0_15_addra[8:0]  ), //i
    .addrb (weightRam_0_15_addrb[8:0]  ), //i
    .dina  (weightRam_0_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_0_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_0 (
    .doutb (weightRam_1_0_doutb[127:0]), //o
    .addra (weightRam_1_0_addra[8:0]  ), //i
    .addrb (weightRam_1_0_addrb[8:0]  ), //i
    .dina  (weightRam_1_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_1 (
    .doutb (weightRam_1_1_doutb[127:0]), //o
    .addra (weightRam_1_1_addra[8:0]  ), //i
    .addrb (weightRam_1_1_addrb[8:0]  ), //i
    .dina  (weightRam_1_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_2 (
    .doutb (weightRam_1_2_doutb[127:0]), //o
    .addra (weightRam_1_2_addra[8:0]  ), //i
    .addrb (weightRam_1_2_addrb[8:0]  ), //i
    .dina  (weightRam_1_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_3 (
    .doutb (weightRam_1_3_doutb[127:0]), //o
    .addra (weightRam_1_3_addra[8:0]  ), //i
    .addrb (weightRam_1_3_addrb[8:0]  ), //i
    .dina  (weightRam_1_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_4 (
    .doutb (weightRam_1_4_doutb[127:0]), //o
    .addra (weightRam_1_4_addra[8:0]  ), //i
    .addrb (weightRam_1_4_addrb[8:0]  ), //i
    .dina  (weightRam_1_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_5 (
    .doutb (weightRam_1_5_doutb[127:0]), //o
    .addra (weightRam_1_5_addra[8:0]  ), //i
    .addrb (weightRam_1_5_addrb[8:0]  ), //i
    .dina  (weightRam_1_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_6 (
    .doutb (weightRam_1_6_doutb[127:0]), //o
    .addra (weightRam_1_6_addra[8:0]  ), //i
    .addrb (weightRam_1_6_addrb[8:0]  ), //i
    .dina  (weightRam_1_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_7 (
    .doutb (weightRam_1_7_doutb[127:0]), //o
    .addra (weightRam_1_7_addra[8:0]  ), //i
    .addrb (weightRam_1_7_addrb[8:0]  ), //i
    .dina  (weightRam_1_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_8 (
    .doutb (weightRam_1_8_doutb[127:0]), //o
    .addra (weightRam_1_8_addra[8:0]  ), //i
    .addrb (weightRam_1_8_addrb[8:0]  ), //i
    .dina  (weightRam_1_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_9 (
    .doutb (weightRam_1_9_doutb[127:0]), //o
    .addra (weightRam_1_9_addra[8:0]  ), //i
    .addrb (weightRam_1_9_addrb[8:0]  ), //i
    .dina  (weightRam_1_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_1_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_1_10 (
    .doutb (weightRam_1_10_doutb[127:0]), //o
    .addra (weightRam_1_10_addra[8:0]  ), //i
    .addrb (weightRam_1_10_addrb[8:0]  ), //i
    .dina  (weightRam_1_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_11 (
    .doutb (weightRam_1_11_doutb[127:0]), //o
    .addra (weightRam_1_11_addra[8:0]  ), //i
    .addrb (weightRam_1_11_addrb[8:0]  ), //i
    .dina  (weightRam_1_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_12 (
    .doutb (weightRam_1_12_doutb[127:0]), //o
    .addra (weightRam_1_12_addra[8:0]  ), //i
    .addrb (weightRam_1_12_addrb[8:0]  ), //i
    .dina  (weightRam_1_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_13 (
    .doutb (weightRam_1_13_doutb[127:0]), //o
    .addra (weightRam_1_13_addra[8:0]  ), //i
    .addrb (weightRam_1_13_addrb[8:0]  ), //i
    .dina  (weightRam_1_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_14 (
    .doutb (weightRam_1_14_doutb[127:0]), //o
    .addra (weightRam_1_14_addra[8:0]  ), //i
    .addrb (weightRam_1_14_addrb[8:0]  ), //i
    .dina  (weightRam_1_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_1_15 (
    .doutb (weightRam_1_15_doutb[127:0]), //o
    .addra (weightRam_1_15_addra[8:0]  ), //i
    .addrb (weightRam_1_15_addrb[8:0]  ), //i
    .dina  (weightRam_1_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_1_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_0 (
    .doutb (weightRam_2_0_doutb[127:0]), //o
    .addra (weightRam_2_0_addra[8:0]  ), //i
    .addrb (weightRam_2_0_addrb[8:0]  ), //i
    .dina  (weightRam_2_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_1 (
    .doutb (weightRam_2_1_doutb[127:0]), //o
    .addra (weightRam_2_1_addra[8:0]  ), //i
    .addrb (weightRam_2_1_addrb[8:0]  ), //i
    .dina  (weightRam_2_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_2 (
    .doutb (weightRam_2_2_doutb[127:0]), //o
    .addra (weightRam_2_2_addra[8:0]  ), //i
    .addrb (weightRam_2_2_addrb[8:0]  ), //i
    .dina  (weightRam_2_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_3 (
    .doutb (weightRam_2_3_doutb[127:0]), //o
    .addra (weightRam_2_3_addra[8:0]  ), //i
    .addrb (weightRam_2_3_addrb[8:0]  ), //i
    .dina  (weightRam_2_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_4 (
    .doutb (weightRam_2_4_doutb[127:0]), //o
    .addra (weightRam_2_4_addra[8:0]  ), //i
    .addrb (weightRam_2_4_addrb[8:0]  ), //i
    .dina  (weightRam_2_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_5 (
    .doutb (weightRam_2_5_doutb[127:0]), //o
    .addra (weightRam_2_5_addra[8:0]  ), //i
    .addrb (weightRam_2_5_addrb[8:0]  ), //i
    .dina  (weightRam_2_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_6 (
    .doutb (weightRam_2_6_doutb[127:0]), //o
    .addra (weightRam_2_6_addra[8:0]  ), //i
    .addrb (weightRam_2_6_addrb[8:0]  ), //i
    .dina  (weightRam_2_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_7 (
    .doutb (weightRam_2_7_doutb[127:0]), //o
    .addra (weightRam_2_7_addra[8:0]  ), //i
    .addrb (weightRam_2_7_addrb[8:0]  ), //i
    .dina  (weightRam_2_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_8 (
    .doutb (weightRam_2_8_doutb[127:0]), //o
    .addra (weightRam_2_8_addra[8:0]  ), //i
    .addrb (weightRam_2_8_addrb[8:0]  ), //i
    .dina  (weightRam_2_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_9 (
    .doutb (weightRam_2_9_doutb[127:0]), //o
    .addra (weightRam_2_9_addra[8:0]  ), //i
    .addrb (weightRam_2_9_addrb[8:0]  ), //i
    .dina  (weightRam_2_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_2_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_2_10 (
    .doutb (weightRam_2_10_doutb[127:0]), //o
    .addra (weightRam_2_10_addra[8:0]  ), //i
    .addrb (weightRam_2_10_addrb[8:0]  ), //i
    .dina  (weightRam_2_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_11 (
    .doutb (weightRam_2_11_doutb[127:0]), //o
    .addra (weightRam_2_11_addra[8:0]  ), //i
    .addrb (weightRam_2_11_addrb[8:0]  ), //i
    .dina  (weightRam_2_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_12 (
    .doutb (weightRam_2_12_doutb[127:0]), //o
    .addra (weightRam_2_12_addra[8:0]  ), //i
    .addrb (weightRam_2_12_addrb[8:0]  ), //i
    .dina  (weightRam_2_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_13 (
    .doutb (weightRam_2_13_doutb[127:0]), //o
    .addra (weightRam_2_13_addra[8:0]  ), //i
    .addrb (weightRam_2_13_addrb[8:0]  ), //i
    .dina  (weightRam_2_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_14 (
    .doutb (weightRam_2_14_doutb[127:0]), //o
    .addra (weightRam_2_14_addra[8:0]  ), //i
    .addrb (weightRam_2_14_addrb[8:0]  ), //i
    .dina  (weightRam_2_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_2_15 (
    .doutb (weightRam_2_15_doutb[127:0]), //o
    .addra (weightRam_2_15_addra[8:0]  ), //i
    .addrb (weightRam_2_15_addrb[8:0]  ), //i
    .dina  (weightRam_2_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_2_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_0 (
    .doutb (weightRam_3_0_doutb[127:0]), //o
    .addra (weightRam_3_0_addra[8:0]  ), //i
    .addrb (weightRam_3_0_addrb[8:0]  ), //i
    .dina  (weightRam_3_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_1 (
    .doutb (weightRam_3_1_doutb[127:0]), //o
    .addra (weightRam_3_1_addra[8:0]  ), //i
    .addrb (weightRam_3_1_addrb[8:0]  ), //i
    .dina  (weightRam_3_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_2 (
    .doutb (weightRam_3_2_doutb[127:0]), //o
    .addra (weightRam_3_2_addra[8:0]  ), //i
    .addrb (weightRam_3_2_addrb[8:0]  ), //i
    .dina  (weightRam_3_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_3 (
    .doutb (weightRam_3_3_doutb[127:0]), //o
    .addra (weightRam_3_3_addra[8:0]  ), //i
    .addrb (weightRam_3_3_addrb[8:0]  ), //i
    .dina  (weightRam_3_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_4 (
    .doutb (weightRam_3_4_doutb[127:0]), //o
    .addra (weightRam_3_4_addra[8:0]  ), //i
    .addrb (weightRam_3_4_addrb[8:0]  ), //i
    .dina  (weightRam_3_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_5 (
    .doutb (weightRam_3_5_doutb[127:0]), //o
    .addra (weightRam_3_5_addra[8:0]  ), //i
    .addrb (weightRam_3_5_addrb[8:0]  ), //i
    .dina  (weightRam_3_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_6 (
    .doutb (weightRam_3_6_doutb[127:0]), //o
    .addra (weightRam_3_6_addra[8:0]  ), //i
    .addrb (weightRam_3_6_addrb[8:0]  ), //i
    .dina  (weightRam_3_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_7 (
    .doutb (weightRam_3_7_doutb[127:0]), //o
    .addra (weightRam_3_7_addra[8:0]  ), //i
    .addrb (weightRam_3_7_addrb[8:0]  ), //i
    .dina  (weightRam_3_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_8 (
    .doutb (weightRam_3_8_doutb[127:0]), //o
    .addra (weightRam_3_8_addra[8:0]  ), //i
    .addrb (weightRam_3_8_addrb[8:0]  ), //i
    .dina  (weightRam_3_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_9 (
    .doutb (weightRam_3_9_doutb[127:0]), //o
    .addra (weightRam_3_9_addra[8:0]  ), //i
    .addrb (weightRam_3_9_addrb[8:0]  ), //i
    .dina  (weightRam_3_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_3_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_3_10 (
    .doutb (weightRam_3_10_doutb[127:0]), //o
    .addra (weightRam_3_10_addra[8:0]  ), //i
    .addrb (weightRam_3_10_addrb[8:0]  ), //i
    .dina  (weightRam_3_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_11 (
    .doutb (weightRam_3_11_doutb[127:0]), //o
    .addra (weightRam_3_11_addra[8:0]  ), //i
    .addrb (weightRam_3_11_addrb[8:0]  ), //i
    .dina  (weightRam_3_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_12 (
    .doutb (weightRam_3_12_doutb[127:0]), //o
    .addra (weightRam_3_12_addra[8:0]  ), //i
    .addrb (weightRam_3_12_addrb[8:0]  ), //i
    .dina  (weightRam_3_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_13 (
    .doutb (weightRam_3_13_doutb[127:0]), //o
    .addra (weightRam_3_13_addra[8:0]  ), //i
    .addrb (weightRam_3_13_addrb[8:0]  ), //i
    .dina  (weightRam_3_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_14 (
    .doutb (weightRam_3_14_doutb[127:0]), //o
    .addra (weightRam_3_14_addra[8:0]  ), //i
    .addrb (weightRam_3_14_addrb[8:0]  ), //i
    .dina  (weightRam_3_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_3_15 (
    .doutb (weightRam_3_15_doutb[127:0]), //o
    .addra (weightRam_3_15_addra[8:0]  ), //i
    .addrb (weightRam_3_15_addrb[8:0]  ), //i
    .dina  (weightRam_3_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_3_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_0 (
    .doutb (weightRam_4_0_doutb[127:0]), //o
    .addra (weightRam_4_0_addra[8:0]  ), //i
    .addrb (weightRam_4_0_addrb[8:0]  ), //i
    .dina  (weightRam_4_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_1 (
    .doutb (weightRam_4_1_doutb[127:0]), //o
    .addra (weightRam_4_1_addra[8:0]  ), //i
    .addrb (weightRam_4_1_addrb[8:0]  ), //i
    .dina  (weightRam_4_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_2 (
    .doutb (weightRam_4_2_doutb[127:0]), //o
    .addra (weightRam_4_2_addra[8:0]  ), //i
    .addrb (weightRam_4_2_addrb[8:0]  ), //i
    .dina  (weightRam_4_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_3 (
    .doutb (weightRam_4_3_doutb[127:0]), //o
    .addra (weightRam_4_3_addra[8:0]  ), //i
    .addrb (weightRam_4_3_addrb[8:0]  ), //i
    .dina  (weightRam_4_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_4 (
    .doutb (weightRam_4_4_doutb[127:0]), //o
    .addra (weightRam_4_4_addra[8:0]  ), //i
    .addrb (weightRam_4_4_addrb[8:0]  ), //i
    .dina  (weightRam_4_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_5 (
    .doutb (weightRam_4_5_doutb[127:0]), //o
    .addra (weightRam_4_5_addra[8:0]  ), //i
    .addrb (weightRam_4_5_addrb[8:0]  ), //i
    .dina  (weightRam_4_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_6 (
    .doutb (weightRam_4_6_doutb[127:0]), //o
    .addra (weightRam_4_6_addra[8:0]  ), //i
    .addrb (weightRam_4_6_addrb[8:0]  ), //i
    .dina  (weightRam_4_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_7 (
    .doutb (weightRam_4_7_doutb[127:0]), //o
    .addra (weightRam_4_7_addra[8:0]  ), //i
    .addrb (weightRam_4_7_addrb[8:0]  ), //i
    .dina  (weightRam_4_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_8 (
    .doutb (weightRam_4_8_doutb[127:0]), //o
    .addra (weightRam_4_8_addra[8:0]  ), //i
    .addrb (weightRam_4_8_addrb[8:0]  ), //i
    .dina  (weightRam_4_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_9 (
    .doutb (weightRam_4_9_doutb[127:0]), //o
    .addra (weightRam_4_9_addra[8:0]  ), //i
    .addrb (weightRam_4_9_addrb[8:0]  ), //i
    .dina  (weightRam_4_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_4_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_4_10 (
    .doutb (weightRam_4_10_doutb[127:0]), //o
    .addra (weightRam_4_10_addra[8:0]  ), //i
    .addrb (weightRam_4_10_addrb[8:0]  ), //i
    .dina  (weightRam_4_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_11 (
    .doutb (weightRam_4_11_doutb[127:0]), //o
    .addra (weightRam_4_11_addra[8:0]  ), //i
    .addrb (weightRam_4_11_addrb[8:0]  ), //i
    .dina  (weightRam_4_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_12 (
    .doutb (weightRam_4_12_doutb[127:0]), //o
    .addra (weightRam_4_12_addra[8:0]  ), //i
    .addrb (weightRam_4_12_addrb[8:0]  ), //i
    .dina  (weightRam_4_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_13 (
    .doutb (weightRam_4_13_doutb[127:0]), //o
    .addra (weightRam_4_13_addra[8:0]  ), //i
    .addrb (weightRam_4_13_addrb[8:0]  ), //i
    .dina  (weightRam_4_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_14 (
    .doutb (weightRam_4_14_doutb[127:0]), //o
    .addra (weightRam_4_14_addra[8:0]  ), //i
    .addrb (weightRam_4_14_addrb[8:0]  ), //i
    .dina  (weightRam_4_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_4_15 (
    .doutb (weightRam_4_15_doutb[127:0]), //o
    .addra (weightRam_4_15_addra[8:0]  ), //i
    .addrb (weightRam_4_15_addrb[8:0]  ), //i
    .dina  (weightRam_4_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_4_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_0 (
    .doutb (weightRam_5_0_doutb[127:0]), //o
    .addra (weightRam_5_0_addra[8:0]  ), //i
    .addrb (weightRam_5_0_addrb[8:0]  ), //i
    .dina  (weightRam_5_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_1 (
    .doutb (weightRam_5_1_doutb[127:0]), //o
    .addra (weightRam_5_1_addra[8:0]  ), //i
    .addrb (weightRam_5_1_addrb[8:0]  ), //i
    .dina  (weightRam_5_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_2 (
    .doutb (weightRam_5_2_doutb[127:0]), //o
    .addra (weightRam_5_2_addra[8:0]  ), //i
    .addrb (weightRam_5_2_addrb[8:0]  ), //i
    .dina  (weightRam_5_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_3 (
    .doutb (weightRam_5_3_doutb[127:0]), //o
    .addra (weightRam_5_3_addra[8:0]  ), //i
    .addrb (weightRam_5_3_addrb[8:0]  ), //i
    .dina  (weightRam_5_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_4 (
    .doutb (weightRam_5_4_doutb[127:0]), //o
    .addra (weightRam_5_4_addra[8:0]  ), //i
    .addrb (weightRam_5_4_addrb[8:0]  ), //i
    .dina  (weightRam_5_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_5 (
    .doutb (weightRam_5_5_doutb[127:0]), //o
    .addra (weightRam_5_5_addra[8:0]  ), //i
    .addrb (weightRam_5_5_addrb[8:0]  ), //i
    .dina  (weightRam_5_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_6 (
    .doutb (weightRam_5_6_doutb[127:0]), //o
    .addra (weightRam_5_6_addra[8:0]  ), //i
    .addrb (weightRam_5_6_addrb[8:0]  ), //i
    .dina  (weightRam_5_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_7 (
    .doutb (weightRam_5_7_doutb[127:0]), //o
    .addra (weightRam_5_7_addra[8:0]  ), //i
    .addrb (weightRam_5_7_addrb[8:0]  ), //i
    .dina  (weightRam_5_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_8 (
    .doutb (weightRam_5_8_doutb[127:0]), //o
    .addra (weightRam_5_8_addra[8:0]  ), //i
    .addrb (weightRam_5_8_addrb[8:0]  ), //i
    .dina  (weightRam_5_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_9 (
    .doutb (weightRam_5_9_doutb[127:0]), //o
    .addra (weightRam_5_9_addra[8:0]  ), //i
    .addrb (weightRam_5_9_addrb[8:0]  ), //i
    .dina  (weightRam_5_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_5_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_5_10 (
    .doutb (weightRam_5_10_doutb[127:0]), //o
    .addra (weightRam_5_10_addra[8:0]  ), //i
    .addrb (weightRam_5_10_addrb[8:0]  ), //i
    .dina  (weightRam_5_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_11 (
    .doutb (weightRam_5_11_doutb[127:0]), //o
    .addra (weightRam_5_11_addra[8:0]  ), //i
    .addrb (weightRam_5_11_addrb[8:0]  ), //i
    .dina  (weightRam_5_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_12 (
    .doutb (weightRam_5_12_doutb[127:0]), //o
    .addra (weightRam_5_12_addra[8:0]  ), //i
    .addrb (weightRam_5_12_addrb[8:0]  ), //i
    .dina  (weightRam_5_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_13 (
    .doutb (weightRam_5_13_doutb[127:0]), //o
    .addra (weightRam_5_13_addra[8:0]  ), //i
    .addrb (weightRam_5_13_addrb[8:0]  ), //i
    .dina  (weightRam_5_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_14 (
    .doutb (weightRam_5_14_doutb[127:0]), //o
    .addra (weightRam_5_14_addra[8:0]  ), //i
    .addrb (weightRam_5_14_addrb[8:0]  ), //i
    .dina  (weightRam_5_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_5_15 (
    .doutb (weightRam_5_15_doutb[127:0]), //o
    .addra (weightRam_5_15_addra[8:0]  ), //i
    .addrb (weightRam_5_15_addrb[8:0]  ), //i
    .dina  (weightRam_5_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_5_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_0 (
    .doutb (weightRam_6_0_doutb[127:0]), //o
    .addra (weightRam_6_0_addra[8:0]  ), //i
    .addrb (weightRam_6_0_addrb[8:0]  ), //i
    .dina  (weightRam_6_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_1 (
    .doutb (weightRam_6_1_doutb[127:0]), //o
    .addra (weightRam_6_1_addra[8:0]  ), //i
    .addrb (weightRam_6_1_addrb[8:0]  ), //i
    .dina  (weightRam_6_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_2 (
    .doutb (weightRam_6_2_doutb[127:0]), //o
    .addra (weightRam_6_2_addra[8:0]  ), //i
    .addrb (weightRam_6_2_addrb[8:0]  ), //i
    .dina  (weightRam_6_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_3 (
    .doutb (weightRam_6_3_doutb[127:0]), //o
    .addra (weightRam_6_3_addra[8:0]  ), //i
    .addrb (weightRam_6_3_addrb[8:0]  ), //i
    .dina  (weightRam_6_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_4 (
    .doutb (weightRam_6_4_doutb[127:0]), //o
    .addra (weightRam_6_4_addra[8:0]  ), //i
    .addrb (weightRam_6_4_addrb[8:0]  ), //i
    .dina  (weightRam_6_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_5 (
    .doutb (weightRam_6_5_doutb[127:0]), //o
    .addra (weightRam_6_5_addra[8:0]  ), //i
    .addrb (weightRam_6_5_addrb[8:0]  ), //i
    .dina  (weightRam_6_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_6 (
    .doutb (weightRam_6_6_doutb[127:0]), //o
    .addra (weightRam_6_6_addra[8:0]  ), //i
    .addrb (weightRam_6_6_addrb[8:0]  ), //i
    .dina  (weightRam_6_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_7 (
    .doutb (weightRam_6_7_doutb[127:0]), //o
    .addra (weightRam_6_7_addra[8:0]  ), //i
    .addrb (weightRam_6_7_addrb[8:0]  ), //i
    .dina  (weightRam_6_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_8 (
    .doutb (weightRam_6_8_doutb[127:0]), //o
    .addra (weightRam_6_8_addra[8:0]  ), //i
    .addrb (weightRam_6_8_addrb[8:0]  ), //i
    .dina  (weightRam_6_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_9 (
    .doutb (weightRam_6_9_doutb[127:0]), //o
    .addra (weightRam_6_9_addra[8:0]  ), //i
    .addrb (weightRam_6_9_addrb[8:0]  ), //i
    .dina  (weightRam_6_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_6_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_6_10 (
    .doutb (weightRam_6_10_doutb[127:0]), //o
    .addra (weightRam_6_10_addra[8:0]  ), //i
    .addrb (weightRam_6_10_addrb[8:0]  ), //i
    .dina  (weightRam_6_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_11 (
    .doutb (weightRam_6_11_doutb[127:0]), //o
    .addra (weightRam_6_11_addra[8:0]  ), //i
    .addrb (weightRam_6_11_addrb[8:0]  ), //i
    .dina  (weightRam_6_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_12 (
    .doutb (weightRam_6_12_doutb[127:0]), //o
    .addra (weightRam_6_12_addra[8:0]  ), //i
    .addrb (weightRam_6_12_addrb[8:0]  ), //i
    .dina  (weightRam_6_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_13 (
    .doutb (weightRam_6_13_doutb[127:0]), //o
    .addra (weightRam_6_13_addra[8:0]  ), //i
    .addrb (weightRam_6_13_addrb[8:0]  ), //i
    .dina  (weightRam_6_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_14 (
    .doutb (weightRam_6_14_doutb[127:0]), //o
    .addra (weightRam_6_14_addra[8:0]  ), //i
    .addrb (weightRam_6_14_addrb[8:0]  ), //i
    .dina  (weightRam_6_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_6_15 (
    .doutb (weightRam_6_15_doutb[127:0]), //o
    .addra (weightRam_6_15_addra[8:0]  ), //i
    .addrb (weightRam_6_15_addrb[8:0]  ), //i
    .dina  (weightRam_6_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_6_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_0 (
    .doutb (weightRam_7_0_doutb[127:0]), //o
    .addra (weightRam_7_0_addra[8:0]  ), //i
    .addrb (weightRam_7_0_addrb[8:0]  ), //i
    .dina  (weightRam_7_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_1 (
    .doutb (weightRam_7_1_doutb[127:0]), //o
    .addra (weightRam_7_1_addra[8:0]  ), //i
    .addrb (weightRam_7_1_addrb[8:0]  ), //i
    .dina  (weightRam_7_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_2 (
    .doutb (weightRam_7_2_doutb[127:0]), //o
    .addra (weightRam_7_2_addra[8:0]  ), //i
    .addrb (weightRam_7_2_addrb[8:0]  ), //i
    .dina  (weightRam_7_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_3 (
    .doutb (weightRam_7_3_doutb[127:0]), //o
    .addra (weightRam_7_3_addra[8:0]  ), //i
    .addrb (weightRam_7_3_addrb[8:0]  ), //i
    .dina  (weightRam_7_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_4 (
    .doutb (weightRam_7_4_doutb[127:0]), //o
    .addra (weightRam_7_4_addra[8:0]  ), //i
    .addrb (weightRam_7_4_addrb[8:0]  ), //i
    .dina  (weightRam_7_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_5 (
    .doutb (weightRam_7_5_doutb[127:0]), //o
    .addra (weightRam_7_5_addra[8:0]  ), //i
    .addrb (weightRam_7_5_addrb[8:0]  ), //i
    .dina  (weightRam_7_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_6 (
    .doutb (weightRam_7_6_doutb[127:0]), //o
    .addra (weightRam_7_6_addra[8:0]  ), //i
    .addrb (weightRam_7_6_addrb[8:0]  ), //i
    .dina  (weightRam_7_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_7 (
    .doutb (weightRam_7_7_doutb[127:0]), //o
    .addra (weightRam_7_7_addra[8:0]  ), //i
    .addrb (weightRam_7_7_addrb[8:0]  ), //i
    .dina  (weightRam_7_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_8 (
    .doutb (weightRam_7_8_doutb[127:0]), //o
    .addra (weightRam_7_8_addra[8:0]  ), //i
    .addrb (weightRam_7_8_addrb[8:0]  ), //i
    .dina  (weightRam_7_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_9 (
    .doutb (weightRam_7_9_doutb[127:0]), //o
    .addra (weightRam_7_9_addra[8:0]  ), //i
    .addrb (weightRam_7_9_addrb[8:0]  ), //i
    .dina  (weightRam_7_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_7_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_7_10 (
    .doutb (weightRam_7_10_doutb[127:0]), //o
    .addra (weightRam_7_10_addra[8:0]  ), //i
    .addrb (weightRam_7_10_addrb[8:0]  ), //i
    .dina  (weightRam_7_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_11 (
    .doutb (weightRam_7_11_doutb[127:0]), //o
    .addra (weightRam_7_11_addra[8:0]  ), //i
    .addrb (weightRam_7_11_addrb[8:0]  ), //i
    .dina  (weightRam_7_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_12 (
    .doutb (weightRam_7_12_doutb[127:0]), //o
    .addra (weightRam_7_12_addra[8:0]  ), //i
    .addrb (weightRam_7_12_addrb[8:0]  ), //i
    .dina  (weightRam_7_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_13 (
    .doutb (weightRam_7_13_doutb[127:0]), //o
    .addra (weightRam_7_13_addra[8:0]  ), //i
    .addrb (weightRam_7_13_addrb[8:0]  ), //i
    .dina  (weightRam_7_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_14 (
    .doutb (weightRam_7_14_doutb[127:0]), //o
    .addra (weightRam_7_14_addra[8:0]  ), //i
    .addrb (weightRam_7_14_addrb[8:0]  ), //i
    .dina  (weightRam_7_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_7_15 (
    .doutb (weightRam_7_15_doutb[127:0]), //o
    .addra (weightRam_7_15_addra[8:0]  ), //i
    .addrb (weightRam_7_15_addrb[8:0]  ), //i
    .dina  (weightRam_7_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_7_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_0 (
    .doutb (weightRam_8_0_doutb[127:0]), //o
    .addra (weightRam_8_0_addra[8:0]  ), //i
    .addrb (weightRam_8_0_addrb[8:0]  ), //i
    .dina  (weightRam_8_0_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_0_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_1 (
    .doutb (weightRam_8_1_doutb[127:0]), //o
    .addra (weightRam_8_1_addra[8:0]  ), //i
    .addrb (weightRam_8_1_addrb[8:0]  ), //i
    .dina  (weightRam_8_1_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_1_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_2 (
    .doutb (weightRam_8_2_doutb[127:0]), //o
    .addra (weightRam_8_2_addra[8:0]  ), //i
    .addrb (weightRam_8_2_addrb[8:0]  ), //i
    .dina  (weightRam_8_2_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_2_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_3 (
    .doutb (weightRam_8_3_doutb[127:0]), //o
    .addra (weightRam_8_3_addra[8:0]  ), //i
    .addrb (weightRam_8_3_addrb[8:0]  ), //i
    .dina  (weightRam_8_3_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_3_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_4 (
    .doutb (weightRam_8_4_doutb[127:0]), //o
    .addra (weightRam_8_4_addra[8:0]  ), //i
    .addrb (weightRam_8_4_addrb[8:0]  ), //i
    .dina  (weightRam_8_4_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_4_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_5 (
    .doutb (weightRam_8_5_doutb[127:0]), //o
    .addra (weightRam_8_5_addra[8:0]  ), //i
    .addrb (weightRam_8_5_addrb[8:0]  ), //i
    .dina  (weightRam_8_5_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_5_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_6 (
    .doutb (weightRam_8_6_doutb[127:0]), //o
    .addra (weightRam_8_6_addra[8:0]  ), //i
    .addrb (weightRam_8_6_addrb[8:0]  ), //i
    .dina  (weightRam_8_6_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_6_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_7 (
    .doutb (weightRam_8_7_doutb[127:0]), //o
    .addra (weightRam_8_7_addra[8:0]  ), //i
    .addrb (weightRam_8_7_addrb[8:0]  ), //i
    .dina  (weightRam_8_7_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_7_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_8 (
    .doutb (weightRam_8_8_doutb[127:0]), //o
    .addra (weightRam_8_8_addra[8:0]  ), //i
    .addrb (weightRam_8_8_addrb[8:0]  ), //i
    .dina  (weightRam_8_8_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_8_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_9 (
    .doutb (weightRam_8_9_doutb[127:0]), //o
    .addra (weightRam_8_9_addra[8:0]  ), //i
    .addrb (weightRam_8_9_addrb[8:0]  ), //i
    .dina  (weightRam_8_9_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (weightRam_8_9_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram weightRam_8_10 (
    .doutb (weightRam_8_10_doutb[127:0]), //o
    .addra (weightRam_8_10_addra[8:0]  ), //i
    .addrb (weightRam_8_10_addrb[8:0]  ), //i
    .dina  (weightRam_8_10_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_10_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_11 (
    .doutb (weightRam_8_11_doutb[127:0]), //o
    .addra (weightRam_8_11_addra[8:0]  ), //i
    .addrb (weightRam_8_11_addrb[8:0]  ), //i
    .dina  (weightRam_8_11_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_11_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_12 (
    .doutb (weightRam_8_12_doutb[127:0]), //o
    .addra (weightRam_8_12_addra[8:0]  ), //i
    .addrb (weightRam_8_12_addrb[8:0]  ), //i
    .dina  (weightRam_8_12_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_12_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_13 (
    .doutb (weightRam_8_13_doutb[127:0]), //o
    .addra (weightRam_8_13_addra[8:0]  ), //i
    .addrb (weightRam_8_13_addrb[8:0]  ), //i
    .dina  (weightRam_8_13_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_13_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_14 (
    .doutb (weightRam_8_14_doutb[127:0]), //o
    .addra (weightRam_8_14_addra[8:0]  ), //i
    .addrb (weightRam_8_14_addrb[8:0]  ), //i
    .dina  (weightRam_8_14_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_14_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram weightRam_8_15 (
    .doutb (weightRam_8_15_doutb[127:0]), //o
    .addra (weightRam_8_15_addra[8:0]  ), //i
    .addrb (weightRam_8_15_addrb[8:0]  ), //i
    .dina  (weightRam_8_15_dina[127:0] ), //i
    .ena   (1'b1                       ), //i
    .enb   (1'b1                       ), //i
    .wea   (weightRam_8_15_wea         ), //i
    .clk   (clk                        )  //i
  );
  sdpram_144 copyBias_ram (
    .doutb (copyBias_ram_doutb[511:0]), //o
    .addra (copyBias_ram_addra[7:0]  ), //i
    .addrb (copyBias_ram_addrb[5:0]  ), //i
    .dina  (copyBias_ram_dina[127:0] ), //i
    .ena   (1'b1                     ), //i
    .enb   (1'b1                     ), //i
    .wea   (copyBias_ram_wea         ), //i
    .clk   (clk                      )  //i
  );
  sdpram_144 copyScale_ram (
    .doutb (copyScale_ram_doutb[511:0]), //o
    .addra (copyScale_ram_addra[7:0]  ), //i
    .addrb (copyScale_ram_addrb[5:0]  ), //i
    .dina  (copyScale_ram_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (copyScale_ram_wea         ), //i
    .clk   (clk                       )  //i
  );
  sdpram_144 copyShift_ram (
    .doutb (copyShift_ram_doutb[511:0]), //o
    .addra (copyShift_ram_addra[7:0]  ), //i
    .addrb (copyShift_ram_addrb[5:0]  ), //i
    .dina  (copyShift_ram_dina[127:0] ), //i
    .ena   (1'b1                      ), //i
    .enb   (1'b1                      ), //i
    .wea   (copyShift_ram_wea         ), //i
    .clk   (clk                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      LoadWeightEnum_IDLE : fsm_currentState_string = "IDLE       ";
      LoadWeightEnum_INIT : fsm_currentState_string = "INIT       ";
      LoadWeightEnum_COPY_WEIGHT : fsm_currentState_string = "COPY_WEIGHT";
      LoadWeightEnum_COPY_BIAS : fsm_currentState_string = "COPY_BIAS  ";
      LoadWeightEnum_COPY_SCALE : fsm_currentState_string = "COPY_SCALE ";
      LoadWeightEnum_COPY_SHIFT : fsm_currentState_string = "COPY_SHIFT ";
      default : fsm_currentState_string = "???????????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      LoadWeightEnum_IDLE : fsm_nextState_string = "IDLE       ";
      LoadWeightEnum_INIT : fsm_nextState_string = "INIT       ";
      LoadWeightEnum_COPY_WEIGHT : fsm_nextState_string = "COPY_WEIGHT";
      LoadWeightEnum_COPY_BIAS : fsm_nextState_string = "COPY_BIAS  ";
      LoadWeightEnum_COPY_SCALE : fsm_nextState_string = "COPY_SCALE ";
      LoadWeightEnum_COPY_SHIFT : fsm_nextState_string = "COPY_SHIFT ";
      default : fsm_nextState_string = "???????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & LoadWeightEnum_IDLE) == LoadWeightEnum_IDLE) : begin
        if(start) begin
          fsm_nextState = LoadWeightEnum_INIT;
        end else begin
          fsm_nextState = LoadWeightEnum_IDLE;
        end
      end
      (((fsm_currentState) & LoadWeightEnum_INIT) == LoadWeightEnum_INIT) : begin
        if(fsm_initEnd) begin
          fsm_nextState = LoadWeightEnum_COPY_WEIGHT;
        end else begin
          fsm_nextState = LoadWeightEnum_INIT;
        end
      end
      (((fsm_currentState) & LoadWeightEnum_COPY_WEIGHT) == LoadWeightEnum_COPY_WEIGHT) : begin
        if(fsm_copyWeightEnd) begin
          fsm_nextState = LoadWeightEnum_COPY_BIAS;
        end else begin
          fsm_nextState = LoadWeightEnum_COPY_WEIGHT;
        end
      end
      (((fsm_currentState) & LoadWeightEnum_COPY_BIAS) == LoadWeightEnum_COPY_BIAS) : begin
        if(fsm_copyBiasEnd) begin
          fsm_nextState = LoadWeightEnum_COPY_SCALE;
        end else begin
          fsm_nextState = LoadWeightEnum_COPY_BIAS;
        end
      end
      (((fsm_currentState) & LoadWeightEnum_COPY_SCALE) == LoadWeightEnum_COPY_SCALE) : begin
        if(fsm_copyScaleEnd) begin
          fsm_nextState = LoadWeightEnum_COPY_SHIFT;
        end else begin
          fsm_nextState = LoadWeightEnum_COPY_SCALE;
        end
      end
      default : begin
        if(fsm_copyShiftEnd) begin
          fsm_nextState = LoadWeightEnum_IDLE;
        end else begin
          fsm_nextState = LoadWeightEnum_COPY_SHIFT;
        end
      end
    endcase
  end

  assign when_WaCounter_l17 = ((fsm_currentState & LoadWeightEnum_INIT) != 6'b000000);
  assign when_WaCounter_l12 = (init_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l12) begin
      init_valid = 1'b1;
    end else begin
      init_valid = 1'b0;
    end
  end

  assign fsm_initEnd = init_valid;
  assign sData_fire = (sData_valid && sData_ready);
  assign when_WaCounter_l17_1 = (((fsm_currentState & LoadWeightEnum_COPY_WEIGHT) != 6'b000000) && sData_fire);
  assign when_WaCounter_l12_1 = (copyWeightCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      copyWeightCnt_valid = 1'b1;
    end else begin
      copyWeightCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l12_2 = (copyWeightTimes_count == 4'b1000);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      copyWeightTimes_valid = 1'b1;
    end else begin
      copyWeightTimes_valid = 1'b0;
    end
  end

  assign sData_fire_1 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_2 = (((fsm_currentState & LoadWeightEnum_COPY_WEIGHT) != 6'b000000) && sData_fire_1);
  assign when_WaCounter_l12_3 = (channelInCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      channelInCnt_valid = 1'b1;
    end else begin
      channelInCnt_valid = 1'b0;
    end
    if(when_Weight_l250) begin
      channelInCnt_valid = 1'b0;
    end
  end

  assign sData_fire_2 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_3 = (((fsm_currentState & LoadWeightEnum_COPY_WEIGHT) != 6'b000000) && sData_fire_2);
  assign when_WaCounter_l12_4 = (computeChannelOut_count == 4'b1111);
  always @(*) begin
    if(when_WaCounter_l12_4) begin
      computeChannelOut_valid = 1'b1;
    end else begin
      computeChannelOut_valid = 1'b0;
    end
    if(when_Weight_l250) begin
      computeChannelOut_valid = 1'b0;
    end
  end

  assign when_WaCounter_l12_5 = (times_count == copyTimes);
  always @(*) begin
    if(when_WaCounter_l12_5) begin
      times_valid = 1'b1;
    end else begin
      times_valid = 1'b0;
    end
    if(when_Weight_l250) begin
      times_valid = 1'b0;
    end
  end

  assign when_WaCounter_l12_6 = (channelOutCnt_count == _zz_when_WaCounter_l12_6);
  always @(*) begin
    if(when_WaCounter_l12_6) begin
      channelOutCnt_valid = 1'b1;
    end else begin
      channelOutCnt_valid = 1'b0;
    end
    if(when_Weight_l250) begin
      channelOutCnt_valid = 1'b0;
    end
  end

  assign when_Weight_l250 = ((fsm_currentState & LoadWeightEnum_IDLE) != 6'b000000);
  assign when_Weight_l256 = (convType == 2'b00);
  always @(*) begin
    if(when_Weight_l256) begin
      fsm_copyWeightEnd = (copyWeightCnt_valid && copyWeightTimes_valid);
    end else begin
      if(when_Weight_l260) begin
        fsm_copyWeightEnd = (channelInCnt_valid && channelOutCnt_valid);
      end else begin
        if(when_Weight_l262) begin
          fsm_copyWeightEnd = copyWeightCnt_valid;
        end else begin
          fsm_copyWeightEnd = 1'b0;
        end
      end
    end
  end

  assign when_Weight_l260 = (convType == 2'b01);
  assign when_Weight_l262 = (convType == 2'b10);
  assign when_Weight_l268 = (((((fsm_currentState & LoadWeightEnum_COPY_WEIGHT) != 6'b000000) || ((fsm_currentState & LoadWeightEnum_COPY_SHIFT) != 6'b000000)) || ((fsm_currentState & LoadWeightEnum_COPY_BIAS) != 6'b000000)) || ((fsm_currentState & LoadWeightEnum_COPY_SCALE) != 6'b000000));
  always @(*) begin
    if(when_Weight_l268) begin
      sData_ready = 1'b1;
    end else begin
      sData_ready = 1'b0;
    end
  end

  assign sData_fire_3 = (sData_valid && sData_ready);
  assign when_Weight_l274 = (sData_fire_3 && ((fsm_currentState & LoadWeightEnum_COPY_WEIGHT) != 6'b000000));
  assign when_Weight_l279 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279) begin
            weav_0_0 = 1'b1;
          end else begin
            weav_0_0 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296) begin
            weav_0_0 = 1'b1;
          end else begin
            weav_0_0 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306) begin
            weav_0_0 = 1'b1;
          end else begin
            weav_0_0 = 1'b0;
          end
        end
        default : begin
          weav_0_0 = 1'b0;
        end
      endcase
    end else begin
      weav_0_0 = 1'b0;
    end
  end

  assign when_Weight_l279_1 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_1) begin
            weav_0_1 = 1'b1;
          end else begin
            weav_0_1 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_1) begin
            weav_0_1 = 1'b1;
          end else begin
            weav_0_1 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_1) begin
            weav_0_1 = 1'b1;
          end else begin
            weav_0_1 = 1'b0;
          end
        end
        default : begin
          weav_0_1 = 1'b0;
        end
      endcase
    end else begin
      weav_0_1 = 1'b0;
    end
  end

  assign when_Weight_l279_2 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_2) begin
            weav_0_2 = 1'b1;
          end else begin
            weav_0_2 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_2) begin
            weav_0_2 = 1'b1;
          end else begin
            weav_0_2 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_2) begin
            weav_0_2 = 1'b1;
          end else begin
            weav_0_2 = 1'b0;
          end
        end
        default : begin
          weav_0_2 = 1'b0;
        end
      endcase
    end else begin
      weav_0_2 = 1'b0;
    end
  end

  assign when_Weight_l279_3 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_3) begin
            weav_0_3 = 1'b1;
          end else begin
            weav_0_3 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_3) begin
            weav_0_3 = 1'b1;
          end else begin
            weav_0_3 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_3) begin
            weav_0_3 = 1'b1;
          end else begin
            weav_0_3 = 1'b0;
          end
        end
        default : begin
          weav_0_3 = 1'b0;
        end
      endcase
    end else begin
      weav_0_3 = 1'b0;
    end
  end

  assign when_Weight_l279_4 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_4) begin
            weav_0_4 = 1'b1;
          end else begin
            weav_0_4 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_4) begin
            weav_0_4 = 1'b1;
          end else begin
            weav_0_4 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_4) begin
            weav_0_4 = 1'b1;
          end else begin
            weav_0_4 = 1'b0;
          end
        end
        default : begin
          weav_0_4 = 1'b0;
        end
      endcase
    end else begin
      weav_0_4 = 1'b0;
    end
  end

  assign when_Weight_l279_5 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_5) begin
            weav_0_5 = 1'b1;
          end else begin
            weav_0_5 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_5) begin
            weav_0_5 = 1'b1;
          end else begin
            weav_0_5 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_5) begin
            weav_0_5 = 1'b1;
          end else begin
            weav_0_5 = 1'b0;
          end
        end
        default : begin
          weav_0_5 = 1'b0;
        end
      endcase
    end else begin
      weav_0_5 = 1'b0;
    end
  end

  assign when_Weight_l279_6 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_6) begin
            weav_0_6 = 1'b1;
          end else begin
            weav_0_6 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_6) begin
            weav_0_6 = 1'b1;
          end else begin
            weav_0_6 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_6) begin
            weav_0_6 = 1'b1;
          end else begin
            weav_0_6 = 1'b0;
          end
        end
        default : begin
          weav_0_6 = 1'b0;
        end
      endcase
    end else begin
      weav_0_6 = 1'b0;
    end
  end

  assign when_Weight_l279_7 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_7) begin
            weav_0_7 = 1'b1;
          end else begin
            weav_0_7 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_7) begin
            weav_0_7 = 1'b1;
          end else begin
            weav_0_7 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_7) begin
            weav_0_7 = 1'b1;
          end else begin
            weav_0_7 = 1'b0;
          end
        end
        default : begin
          weav_0_7 = 1'b0;
        end
      endcase
    end else begin
      weav_0_7 = 1'b0;
    end
  end

  assign when_Weight_l279_8 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_8) begin
            weav_0_8 = 1'b1;
          end else begin
            weav_0_8 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_8) begin
            weav_0_8 = 1'b1;
          end else begin
            weav_0_8 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_8) begin
            weav_0_8 = 1'b1;
          end else begin
            weav_0_8 = 1'b0;
          end
        end
        default : begin
          weav_0_8 = 1'b0;
        end
      endcase
    end else begin
      weav_0_8 = 1'b0;
    end
  end

  assign when_Weight_l279_9 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_9) begin
            weav_0_9 = 1'b1;
          end else begin
            weav_0_9 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_9) begin
            weav_0_9 = 1'b1;
          end else begin
            weav_0_9 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_9) begin
            weav_0_9 = 1'b1;
          end else begin
            weav_0_9 = 1'b0;
          end
        end
        default : begin
          weav_0_9 = 1'b0;
        end
      endcase
    end else begin
      weav_0_9 = 1'b0;
    end
  end

  assign when_Weight_l279_10 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_10) begin
            weav_0_10 = 1'b1;
          end else begin
            weav_0_10 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_10) begin
            weav_0_10 = 1'b1;
          end else begin
            weav_0_10 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_10) begin
            weav_0_10 = 1'b1;
          end else begin
            weav_0_10 = 1'b0;
          end
        end
        default : begin
          weav_0_10 = 1'b0;
        end
      endcase
    end else begin
      weav_0_10 = 1'b0;
    end
  end

  assign when_Weight_l279_11 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_11) begin
            weav_0_11 = 1'b1;
          end else begin
            weav_0_11 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_11) begin
            weav_0_11 = 1'b1;
          end else begin
            weav_0_11 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_11) begin
            weav_0_11 = 1'b1;
          end else begin
            weav_0_11 = 1'b0;
          end
        end
        default : begin
          weav_0_11 = 1'b0;
        end
      endcase
    end else begin
      weav_0_11 = 1'b0;
    end
  end

  assign when_Weight_l279_12 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_12) begin
            weav_0_12 = 1'b1;
          end else begin
            weav_0_12 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_12) begin
            weav_0_12 = 1'b1;
          end else begin
            weav_0_12 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_12) begin
            weav_0_12 = 1'b1;
          end else begin
            weav_0_12 = 1'b0;
          end
        end
        default : begin
          weav_0_12 = 1'b0;
        end
      endcase
    end else begin
      weav_0_12 = 1'b0;
    end
  end

  assign when_Weight_l279_13 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_13) begin
            weav_0_13 = 1'b1;
          end else begin
            weav_0_13 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_13) begin
            weav_0_13 = 1'b1;
          end else begin
            weav_0_13 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_13) begin
            weav_0_13 = 1'b1;
          end else begin
            weav_0_13 = 1'b0;
          end
        end
        default : begin
          weav_0_13 = 1'b0;
        end
      endcase
    end else begin
      weav_0_13 = 1'b0;
    end
  end

  assign when_Weight_l279_14 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_14) begin
            weav_0_14 = 1'b1;
          end else begin
            weav_0_14 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_14) begin
            weav_0_14 = 1'b1;
          end else begin
            weav_0_14 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_14) begin
            weav_0_14 = 1'b1;
          end else begin
            weav_0_14 = 1'b0;
          end
        end
        default : begin
          weav_0_14 = 1'b0;
        end
      endcase
    end else begin
      weav_0_14 = 1'b0;
    end
  end

  assign when_Weight_l279_15 = ((copyWeightTimes_count == 4'b0000) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_15) begin
            weav_0_15 = 1'b1;
          end else begin
            weav_0_15 = 1'b0;
          end
        end
        2'b10 : begin
          if(when_Weight_l296_15) begin
            weav_0_15 = 1'b1;
          end else begin
            weav_0_15 = 1'b0;
          end
        end
        2'b01 : begin
          if(when_Weight_l306_15) begin
            weav_0_15 = 1'b1;
          end else begin
            weav_0_15 = 1'b0;
          end
        end
        default : begin
          weav_0_15 = 1'b0;
        end
      endcase
    end else begin
      weav_0_15 = 1'b0;
    end
  end

  assign when_Weight_l279_16 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_16) begin
            weav_1_0 = 1'b1;
          end else begin
            weav_1_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_16) begin
            weav_1_0 = 1'b1;
          end else begin
            weav_1_0 = 1'b0;
          end
        end
        default : begin
          weav_1_0 = 1'b0;
        end
      endcase
    end else begin
      weav_1_0 = 1'b0;
    end
  end

  assign when_Weight_l279_17 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_17) begin
            weav_1_1 = 1'b1;
          end else begin
            weav_1_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_17) begin
            weav_1_1 = 1'b1;
          end else begin
            weav_1_1 = 1'b0;
          end
        end
        default : begin
          weav_1_1 = 1'b0;
        end
      endcase
    end else begin
      weav_1_1 = 1'b0;
    end
  end

  assign when_Weight_l279_18 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_18) begin
            weav_1_2 = 1'b1;
          end else begin
            weav_1_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_18) begin
            weav_1_2 = 1'b1;
          end else begin
            weav_1_2 = 1'b0;
          end
        end
        default : begin
          weav_1_2 = 1'b0;
        end
      endcase
    end else begin
      weav_1_2 = 1'b0;
    end
  end

  assign when_Weight_l279_19 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_19) begin
            weav_1_3 = 1'b1;
          end else begin
            weav_1_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_19) begin
            weav_1_3 = 1'b1;
          end else begin
            weav_1_3 = 1'b0;
          end
        end
        default : begin
          weav_1_3 = 1'b0;
        end
      endcase
    end else begin
      weav_1_3 = 1'b0;
    end
  end

  assign when_Weight_l279_20 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_20) begin
            weav_1_4 = 1'b1;
          end else begin
            weav_1_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_20) begin
            weav_1_4 = 1'b1;
          end else begin
            weav_1_4 = 1'b0;
          end
        end
        default : begin
          weav_1_4 = 1'b0;
        end
      endcase
    end else begin
      weav_1_4 = 1'b0;
    end
  end

  assign when_Weight_l279_21 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_21) begin
            weav_1_5 = 1'b1;
          end else begin
            weav_1_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_21) begin
            weav_1_5 = 1'b1;
          end else begin
            weav_1_5 = 1'b0;
          end
        end
        default : begin
          weav_1_5 = 1'b0;
        end
      endcase
    end else begin
      weav_1_5 = 1'b0;
    end
  end

  assign when_Weight_l279_22 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_22) begin
            weav_1_6 = 1'b1;
          end else begin
            weav_1_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_22) begin
            weav_1_6 = 1'b1;
          end else begin
            weav_1_6 = 1'b0;
          end
        end
        default : begin
          weav_1_6 = 1'b0;
        end
      endcase
    end else begin
      weav_1_6 = 1'b0;
    end
  end

  assign when_Weight_l279_23 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_23) begin
            weav_1_7 = 1'b1;
          end else begin
            weav_1_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_23) begin
            weav_1_7 = 1'b1;
          end else begin
            weav_1_7 = 1'b0;
          end
        end
        default : begin
          weav_1_7 = 1'b0;
        end
      endcase
    end else begin
      weav_1_7 = 1'b0;
    end
  end

  assign when_Weight_l279_24 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_24) begin
            weav_1_8 = 1'b1;
          end else begin
            weav_1_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_24) begin
            weav_1_8 = 1'b1;
          end else begin
            weav_1_8 = 1'b0;
          end
        end
        default : begin
          weav_1_8 = 1'b0;
        end
      endcase
    end else begin
      weav_1_8 = 1'b0;
    end
  end

  assign when_Weight_l279_25 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_25) begin
            weav_1_9 = 1'b1;
          end else begin
            weav_1_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_25) begin
            weav_1_9 = 1'b1;
          end else begin
            weav_1_9 = 1'b0;
          end
        end
        default : begin
          weav_1_9 = 1'b0;
        end
      endcase
    end else begin
      weav_1_9 = 1'b0;
    end
  end

  assign when_Weight_l279_26 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_26) begin
            weav_1_10 = 1'b1;
          end else begin
            weav_1_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_26) begin
            weav_1_10 = 1'b1;
          end else begin
            weav_1_10 = 1'b0;
          end
        end
        default : begin
          weav_1_10 = 1'b0;
        end
      endcase
    end else begin
      weav_1_10 = 1'b0;
    end
  end

  assign when_Weight_l279_27 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_27) begin
            weav_1_11 = 1'b1;
          end else begin
            weav_1_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_27) begin
            weav_1_11 = 1'b1;
          end else begin
            weav_1_11 = 1'b0;
          end
        end
        default : begin
          weav_1_11 = 1'b0;
        end
      endcase
    end else begin
      weav_1_11 = 1'b0;
    end
  end

  assign when_Weight_l279_28 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_28) begin
            weav_1_12 = 1'b1;
          end else begin
            weav_1_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_28) begin
            weav_1_12 = 1'b1;
          end else begin
            weav_1_12 = 1'b0;
          end
        end
        default : begin
          weav_1_12 = 1'b0;
        end
      endcase
    end else begin
      weav_1_12 = 1'b0;
    end
  end

  assign when_Weight_l279_29 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_29) begin
            weav_1_13 = 1'b1;
          end else begin
            weav_1_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_29) begin
            weav_1_13 = 1'b1;
          end else begin
            weav_1_13 = 1'b0;
          end
        end
        default : begin
          weav_1_13 = 1'b0;
        end
      endcase
    end else begin
      weav_1_13 = 1'b0;
    end
  end

  assign when_Weight_l279_30 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_30) begin
            weav_1_14 = 1'b1;
          end else begin
            weav_1_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_30) begin
            weav_1_14 = 1'b1;
          end else begin
            weav_1_14 = 1'b0;
          end
        end
        default : begin
          weav_1_14 = 1'b0;
        end
      endcase
    end else begin
      weav_1_14 = 1'b0;
    end
  end

  assign when_Weight_l279_31 = ((copyWeightTimes_count == 4'b0001) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_31) begin
            weav_1_15 = 1'b1;
          end else begin
            weav_1_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_1_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_31) begin
            weav_1_15 = 1'b1;
          end else begin
            weav_1_15 = 1'b0;
          end
        end
        default : begin
          weav_1_15 = 1'b0;
        end
      endcase
    end else begin
      weav_1_15 = 1'b0;
    end
  end

  assign when_Weight_l279_32 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_32) begin
            weav_2_0 = 1'b1;
          end else begin
            weav_2_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_32) begin
            weav_2_0 = 1'b1;
          end else begin
            weav_2_0 = 1'b0;
          end
        end
        default : begin
          weav_2_0 = 1'b0;
        end
      endcase
    end else begin
      weav_2_0 = 1'b0;
    end
  end

  assign when_Weight_l279_33 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_33) begin
            weav_2_1 = 1'b1;
          end else begin
            weav_2_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_33) begin
            weav_2_1 = 1'b1;
          end else begin
            weav_2_1 = 1'b0;
          end
        end
        default : begin
          weav_2_1 = 1'b0;
        end
      endcase
    end else begin
      weav_2_1 = 1'b0;
    end
  end

  assign when_Weight_l279_34 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_34) begin
            weav_2_2 = 1'b1;
          end else begin
            weav_2_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_34) begin
            weav_2_2 = 1'b1;
          end else begin
            weav_2_2 = 1'b0;
          end
        end
        default : begin
          weav_2_2 = 1'b0;
        end
      endcase
    end else begin
      weav_2_2 = 1'b0;
    end
  end

  assign when_Weight_l279_35 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_35) begin
            weav_2_3 = 1'b1;
          end else begin
            weav_2_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_35) begin
            weav_2_3 = 1'b1;
          end else begin
            weav_2_3 = 1'b0;
          end
        end
        default : begin
          weav_2_3 = 1'b0;
        end
      endcase
    end else begin
      weav_2_3 = 1'b0;
    end
  end

  assign when_Weight_l279_36 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_36) begin
            weav_2_4 = 1'b1;
          end else begin
            weav_2_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_36) begin
            weav_2_4 = 1'b1;
          end else begin
            weav_2_4 = 1'b0;
          end
        end
        default : begin
          weav_2_4 = 1'b0;
        end
      endcase
    end else begin
      weav_2_4 = 1'b0;
    end
  end

  assign when_Weight_l279_37 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_37) begin
            weav_2_5 = 1'b1;
          end else begin
            weav_2_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_37) begin
            weav_2_5 = 1'b1;
          end else begin
            weav_2_5 = 1'b0;
          end
        end
        default : begin
          weav_2_5 = 1'b0;
        end
      endcase
    end else begin
      weav_2_5 = 1'b0;
    end
  end

  assign when_Weight_l279_38 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_38) begin
            weav_2_6 = 1'b1;
          end else begin
            weav_2_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_38) begin
            weav_2_6 = 1'b1;
          end else begin
            weav_2_6 = 1'b0;
          end
        end
        default : begin
          weav_2_6 = 1'b0;
        end
      endcase
    end else begin
      weav_2_6 = 1'b0;
    end
  end

  assign when_Weight_l279_39 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_39) begin
            weav_2_7 = 1'b1;
          end else begin
            weav_2_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_39) begin
            weav_2_7 = 1'b1;
          end else begin
            weav_2_7 = 1'b0;
          end
        end
        default : begin
          weav_2_7 = 1'b0;
        end
      endcase
    end else begin
      weav_2_7 = 1'b0;
    end
  end

  assign when_Weight_l279_40 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_40) begin
            weav_2_8 = 1'b1;
          end else begin
            weav_2_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_40) begin
            weav_2_8 = 1'b1;
          end else begin
            weav_2_8 = 1'b0;
          end
        end
        default : begin
          weav_2_8 = 1'b0;
        end
      endcase
    end else begin
      weav_2_8 = 1'b0;
    end
  end

  assign when_Weight_l279_41 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_41) begin
            weav_2_9 = 1'b1;
          end else begin
            weav_2_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_41) begin
            weav_2_9 = 1'b1;
          end else begin
            weav_2_9 = 1'b0;
          end
        end
        default : begin
          weav_2_9 = 1'b0;
        end
      endcase
    end else begin
      weav_2_9 = 1'b0;
    end
  end

  assign when_Weight_l279_42 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_42) begin
            weav_2_10 = 1'b1;
          end else begin
            weav_2_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_42) begin
            weav_2_10 = 1'b1;
          end else begin
            weav_2_10 = 1'b0;
          end
        end
        default : begin
          weav_2_10 = 1'b0;
        end
      endcase
    end else begin
      weav_2_10 = 1'b0;
    end
  end

  assign when_Weight_l279_43 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_43) begin
            weav_2_11 = 1'b1;
          end else begin
            weav_2_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_43) begin
            weav_2_11 = 1'b1;
          end else begin
            weav_2_11 = 1'b0;
          end
        end
        default : begin
          weav_2_11 = 1'b0;
        end
      endcase
    end else begin
      weav_2_11 = 1'b0;
    end
  end

  assign when_Weight_l279_44 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_44) begin
            weav_2_12 = 1'b1;
          end else begin
            weav_2_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_44) begin
            weav_2_12 = 1'b1;
          end else begin
            weav_2_12 = 1'b0;
          end
        end
        default : begin
          weav_2_12 = 1'b0;
        end
      endcase
    end else begin
      weav_2_12 = 1'b0;
    end
  end

  assign when_Weight_l279_45 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_45) begin
            weav_2_13 = 1'b1;
          end else begin
            weav_2_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_45) begin
            weav_2_13 = 1'b1;
          end else begin
            weav_2_13 = 1'b0;
          end
        end
        default : begin
          weav_2_13 = 1'b0;
        end
      endcase
    end else begin
      weav_2_13 = 1'b0;
    end
  end

  assign when_Weight_l279_46 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_46) begin
            weav_2_14 = 1'b1;
          end else begin
            weav_2_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_46) begin
            weav_2_14 = 1'b1;
          end else begin
            weav_2_14 = 1'b0;
          end
        end
        default : begin
          weav_2_14 = 1'b0;
        end
      endcase
    end else begin
      weav_2_14 = 1'b0;
    end
  end

  assign when_Weight_l279_47 = ((copyWeightTimes_count == 4'b0010) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_47) begin
            weav_2_15 = 1'b1;
          end else begin
            weav_2_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_2_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_47) begin
            weav_2_15 = 1'b1;
          end else begin
            weav_2_15 = 1'b0;
          end
        end
        default : begin
          weav_2_15 = 1'b0;
        end
      endcase
    end else begin
      weav_2_15 = 1'b0;
    end
  end

  assign when_Weight_l279_48 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_48) begin
            weav_3_0 = 1'b1;
          end else begin
            weav_3_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_48) begin
            weav_3_0 = 1'b1;
          end else begin
            weav_3_0 = 1'b0;
          end
        end
        default : begin
          weav_3_0 = 1'b0;
        end
      endcase
    end else begin
      weav_3_0 = 1'b0;
    end
  end

  assign when_Weight_l279_49 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_49) begin
            weav_3_1 = 1'b1;
          end else begin
            weav_3_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_49) begin
            weav_3_1 = 1'b1;
          end else begin
            weav_3_1 = 1'b0;
          end
        end
        default : begin
          weav_3_1 = 1'b0;
        end
      endcase
    end else begin
      weav_3_1 = 1'b0;
    end
  end

  assign when_Weight_l279_50 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_50) begin
            weav_3_2 = 1'b1;
          end else begin
            weav_3_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_50) begin
            weav_3_2 = 1'b1;
          end else begin
            weav_3_2 = 1'b0;
          end
        end
        default : begin
          weav_3_2 = 1'b0;
        end
      endcase
    end else begin
      weav_3_2 = 1'b0;
    end
  end

  assign when_Weight_l279_51 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_51) begin
            weav_3_3 = 1'b1;
          end else begin
            weav_3_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_51) begin
            weav_3_3 = 1'b1;
          end else begin
            weav_3_3 = 1'b0;
          end
        end
        default : begin
          weav_3_3 = 1'b0;
        end
      endcase
    end else begin
      weav_3_3 = 1'b0;
    end
  end

  assign when_Weight_l279_52 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_52) begin
            weav_3_4 = 1'b1;
          end else begin
            weav_3_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_52) begin
            weav_3_4 = 1'b1;
          end else begin
            weav_3_4 = 1'b0;
          end
        end
        default : begin
          weav_3_4 = 1'b0;
        end
      endcase
    end else begin
      weav_3_4 = 1'b0;
    end
  end

  assign when_Weight_l279_53 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_53) begin
            weav_3_5 = 1'b1;
          end else begin
            weav_3_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_53) begin
            weav_3_5 = 1'b1;
          end else begin
            weav_3_5 = 1'b0;
          end
        end
        default : begin
          weav_3_5 = 1'b0;
        end
      endcase
    end else begin
      weav_3_5 = 1'b0;
    end
  end

  assign when_Weight_l279_54 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_54) begin
            weav_3_6 = 1'b1;
          end else begin
            weav_3_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_54) begin
            weav_3_6 = 1'b1;
          end else begin
            weav_3_6 = 1'b0;
          end
        end
        default : begin
          weav_3_6 = 1'b0;
        end
      endcase
    end else begin
      weav_3_6 = 1'b0;
    end
  end

  assign when_Weight_l279_55 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_55) begin
            weav_3_7 = 1'b1;
          end else begin
            weav_3_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_55) begin
            weav_3_7 = 1'b1;
          end else begin
            weav_3_7 = 1'b0;
          end
        end
        default : begin
          weav_3_7 = 1'b0;
        end
      endcase
    end else begin
      weav_3_7 = 1'b0;
    end
  end

  assign when_Weight_l279_56 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_56) begin
            weav_3_8 = 1'b1;
          end else begin
            weav_3_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_56) begin
            weav_3_8 = 1'b1;
          end else begin
            weav_3_8 = 1'b0;
          end
        end
        default : begin
          weav_3_8 = 1'b0;
        end
      endcase
    end else begin
      weav_3_8 = 1'b0;
    end
  end

  assign when_Weight_l279_57 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_57) begin
            weav_3_9 = 1'b1;
          end else begin
            weav_3_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_57) begin
            weav_3_9 = 1'b1;
          end else begin
            weav_3_9 = 1'b0;
          end
        end
        default : begin
          weav_3_9 = 1'b0;
        end
      endcase
    end else begin
      weav_3_9 = 1'b0;
    end
  end

  assign when_Weight_l279_58 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_58) begin
            weav_3_10 = 1'b1;
          end else begin
            weav_3_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_58) begin
            weav_3_10 = 1'b1;
          end else begin
            weav_3_10 = 1'b0;
          end
        end
        default : begin
          weav_3_10 = 1'b0;
        end
      endcase
    end else begin
      weav_3_10 = 1'b0;
    end
  end

  assign when_Weight_l279_59 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_59) begin
            weav_3_11 = 1'b1;
          end else begin
            weav_3_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_59) begin
            weav_3_11 = 1'b1;
          end else begin
            weav_3_11 = 1'b0;
          end
        end
        default : begin
          weav_3_11 = 1'b0;
        end
      endcase
    end else begin
      weav_3_11 = 1'b0;
    end
  end

  assign when_Weight_l279_60 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_60) begin
            weav_3_12 = 1'b1;
          end else begin
            weav_3_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_60) begin
            weav_3_12 = 1'b1;
          end else begin
            weav_3_12 = 1'b0;
          end
        end
        default : begin
          weav_3_12 = 1'b0;
        end
      endcase
    end else begin
      weav_3_12 = 1'b0;
    end
  end

  assign when_Weight_l279_61 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_61) begin
            weav_3_13 = 1'b1;
          end else begin
            weav_3_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_61) begin
            weav_3_13 = 1'b1;
          end else begin
            weav_3_13 = 1'b0;
          end
        end
        default : begin
          weav_3_13 = 1'b0;
        end
      endcase
    end else begin
      weav_3_13 = 1'b0;
    end
  end

  assign when_Weight_l279_62 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_62) begin
            weav_3_14 = 1'b1;
          end else begin
            weav_3_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_62) begin
            weav_3_14 = 1'b1;
          end else begin
            weav_3_14 = 1'b0;
          end
        end
        default : begin
          weav_3_14 = 1'b0;
        end
      endcase
    end else begin
      weav_3_14 = 1'b0;
    end
  end

  assign when_Weight_l279_63 = ((copyWeightTimes_count == 4'b0011) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_63) begin
            weav_3_15 = 1'b1;
          end else begin
            weav_3_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_3_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_63) begin
            weav_3_15 = 1'b1;
          end else begin
            weav_3_15 = 1'b0;
          end
        end
        default : begin
          weav_3_15 = 1'b0;
        end
      endcase
    end else begin
      weav_3_15 = 1'b0;
    end
  end

  assign when_Weight_l279_64 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_64) begin
            weav_4_0 = 1'b1;
          end else begin
            weav_4_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_64) begin
            weav_4_0 = 1'b1;
          end else begin
            weav_4_0 = 1'b0;
          end
        end
        default : begin
          weav_4_0 = 1'b0;
        end
      endcase
    end else begin
      weav_4_0 = 1'b0;
    end
  end

  assign when_Weight_l279_65 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_65) begin
            weav_4_1 = 1'b1;
          end else begin
            weav_4_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_65) begin
            weav_4_1 = 1'b1;
          end else begin
            weav_4_1 = 1'b0;
          end
        end
        default : begin
          weav_4_1 = 1'b0;
        end
      endcase
    end else begin
      weav_4_1 = 1'b0;
    end
  end

  assign when_Weight_l279_66 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_66) begin
            weav_4_2 = 1'b1;
          end else begin
            weav_4_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_66) begin
            weav_4_2 = 1'b1;
          end else begin
            weav_4_2 = 1'b0;
          end
        end
        default : begin
          weav_4_2 = 1'b0;
        end
      endcase
    end else begin
      weav_4_2 = 1'b0;
    end
  end

  assign when_Weight_l279_67 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_67) begin
            weav_4_3 = 1'b1;
          end else begin
            weav_4_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_67) begin
            weav_4_3 = 1'b1;
          end else begin
            weav_4_3 = 1'b0;
          end
        end
        default : begin
          weav_4_3 = 1'b0;
        end
      endcase
    end else begin
      weav_4_3 = 1'b0;
    end
  end

  assign when_Weight_l279_68 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_68) begin
            weav_4_4 = 1'b1;
          end else begin
            weav_4_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_68) begin
            weav_4_4 = 1'b1;
          end else begin
            weav_4_4 = 1'b0;
          end
        end
        default : begin
          weav_4_4 = 1'b0;
        end
      endcase
    end else begin
      weav_4_4 = 1'b0;
    end
  end

  assign when_Weight_l279_69 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_69) begin
            weav_4_5 = 1'b1;
          end else begin
            weav_4_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_69) begin
            weav_4_5 = 1'b1;
          end else begin
            weav_4_5 = 1'b0;
          end
        end
        default : begin
          weav_4_5 = 1'b0;
        end
      endcase
    end else begin
      weav_4_5 = 1'b0;
    end
  end

  assign when_Weight_l279_70 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_70) begin
            weav_4_6 = 1'b1;
          end else begin
            weav_4_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_70) begin
            weav_4_6 = 1'b1;
          end else begin
            weav_4_6 = 1'b0;
          end
        end
        default : begin
          weav_4_6 = 1'b0;
        end
      endcase
    end else begin
      weav_4_6 = 1'b0;
    end
  end

  assign when_Weight_l279_71 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_71) begin
            weav_4_7 = 1'b1;
          end else begin
            weav_4_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_71) begin
            weav_4_7 = 1'b1;
          end else begin
            weav_4_7 = 1'b0;
          end
        end
        default : begin
          weav_4_7 = 1'b0;
        end
      endcase
    end else begin
      weav_4_7 = 1'b0;
    end
  end

  assign when_Weight_l279_72 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_72) begin
            weav_4_8 = 1'b1;
          end else begin
            weav_4_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_72) begin
            weav_4_8 = 1'b1;
          end else begin
            weav_4_8 = 1'b0;
          end
        end
        default : begin
          weav_4_8 = 1'b0;
        end
      endcase
    end else begin
      weav_4_8 = 1'b0;
    end
  end

  assign when_Weight_l279_73 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_73) begin
            weav_4_9 = 1'b1;
          end else begin
            weav_4_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_73) begin
            weav_4_9 = 1'b1;
          end else begin
            weav_4_9 = 1'b0;
          end
        end
        default : begin
          weav_4_9 = 1'b0;
        end
      endcase
    end else begin
      weav_4_9 = 1'b0;
    end
  end

  assign when_Weight_l279_74 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_74) begin
            weav_4_10 = 1'b1;
          end else begin
            weav_4_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_74) begin
            weav_4_10 = 1'b1;
          end else begin
            weav_4_10 = 1'b0;
          end
        end
        default : begin
          weav_4_10 = 1'b0;
        end
      endcase
    end else begin
      weav_4_10 = 1'b0;
    end
  end

  assign when_Weight_l279_75 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_75) begin
            weav_4_11 = 1'b1;
          end else begin
            weav_4_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_75) begin
            weav_4_11 = 1'b1;
          end else begin
            weav_4_11 = 1'b0;
          end
        end
        default : begin
          weav_4_11 = 1'b0;
        end
      endcase
    end else begin
      weav_4_11 = 1'b0;
    end
  end

  assign when_Weight_l279_76 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_76) begin
            weav_4_12 = 1'b1;
          end else begin
            weav_4_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_76) begin
            weav_4_12 = 1'b1;
          end else begin
            weav_4_12 = 1'b0;
          end
        end
        default : begin
          weav_4_12 = 1'b0;
        end
      endcase
    end else begin
      weav_4_12 = 1'b0;
    end
  end

  assign when_Weight_l279_77 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_77) begin
            weav_4_13 = 1'b1;
          end else begin
            weav_4_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_77) begin
            weav_4_13 = 1'b1;
          end else begin
            weav_4_13 = 1'b0;
          end
        end
        default : begin
          weav_4_13 = 1'b0;
        end
      endcase
    end else begin
      weav_4_13 = 1'b0;
    end
  end

  assign when_Weight_l279_78 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_78) begin
            weav_4_14 = 1'b1;
          end else begin
            weav_4_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_78) begin
            weav_4_14 = 1'b1;
          end else begin
            weav_4_14 = 1'b0;
          end
        end
        default : begin
          weav_4_14 = 1'b0;
        end
      endcase
    end else begin
      weav_4_14 = 1'b0;
    end
  end

  assign when_Weight_l279_79 = ((copyWeightTimes_count == 4'b0100) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_79) begin
            weav_4_15 = 1'b1;
          end else begin
            weav_4_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_4_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_79) begin
            weav_4_15 = 1'b1;
          end else begin
            weav_4_15 = 1'b0;
          end
        end
        default : begin
          weav_4_15 = 1'b0;
        end
      endcase
    end else begin
      weav_4_15 = 1'b0;
    end
  end

  assign when_Weight_l279_80 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_80) begin
            weav_5_0 = 1'b1;
          end else begin
            weav_5_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_80) begin
            weav_5_0 = 1'b1;
          end else begin
            weav_5_0 = 1'b0;
          end
        end
        default : begin
          weav_5_0 = 1'b0;
        end
      endcase
    end else begin
      weav_5_0 = 1'b0;
    end
  end

  assign when_Weight_l279_81 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_81) begin
            weav_5_1 = 1'b1;
          end else begin
            weav_5_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_81) begin
            weav_5_1 = 1'b1;
          end else begin
            weav_5_1 = 1'b0;
          end
        end
        default : begin
          weav_5_1 = 1'b0;
        end
      endcase
    end else begin
      weav_5_1 = 1'b0;
    end
  end

  assign when_Weight_l279_82 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_82) begin
            weav_5_2 = 1'b1;
          end else begin
            weav_5_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_82) begin
            weav_5_2 = 1'b1;
          end else begin
            weav_5_2 = 1'b0;
          end
        end
        default : begin
          weav_5_2 = 1'b0;
        end
      endcase
    end else begin
      weav_5_2 = 1'b0;
    end
  end

  assign when_Weight_l279_83 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_83) begin
            weav_5_3 = 1'b1;
          end else begin
            weav_5_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_83) begin
            weav_5_3 = 1'b1;
          end else begin
            weav_5_3 = 1'b0;
          end
        end
        default : begin
          weav_5_3 = 1'b0;
        end
      endcase
    end else begin
      weav_5_3 = 1'b0;
    end
  end

  assign when_Weight_l279_84 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_84) begin
            weav_5_4 = 1'b1;
          end else begin
            weav_5_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_84) begin
            weav_5_4 = 1'b1;
          end else begin
            weav_5_4 = 1'b0;
          end
        end
        default : begin
          weav_5_4 = 1'b0;
        end
      endcase
    end else begin
      weav_5_4 = 1'b0;
    end
  end

  assign when_Weight_l279_85 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_85) begin
            weav_5_5 = 1'b1;
          end else begin
            weav_5_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_85) begin
            weav_5_5 = 1'b1;
          end else begin
            weav_5_5 = 1'b0;
          end
        end
        default : begin
          weav_5_5 = 1'b0;
        end
      endcase
    end else begin
      weav_5_5 = 1'b0;
    end
  end

  assign when_Weight_l279_86 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_86) begin
            weav_5_6 = 1'b1;
          end else begin
            weav_5_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_86) begin
            weav_5_6 = 1'b1;
          end else begin
            weav_5_6 = 1'b0;
          end
        end
        default : begin
          weav_5_6 = 1'b0;
        end
      endcase
    end else begin
      weav_5_6 = 1'b0;
    end
  end

  assign when_Weight_l279_87 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_87) begin
            weav_5_7 = 1'b1;
          end else begin
            weav_5_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_87) begin
            weav_5_7 = 1'b1;
          end else begin
            weav_5_7 = 1'b0;
          end
        end
        default : begin
          weav_5_7 = 1'b0;
        end
      endcase
    end else begin
      weav_5_7 = 1'b0;
    end
  end

  assign when_Weight_l279_88 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_88) begin
            weav_5_8 = 1'b1;
          end else begin
            weav_5_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_88) begin
            weav_5_8 = 1'b1;
          end else begin
            weav_5_8 = 1'b0;
          end
        end
        default : begin
          weav_5_8 = 1'b0;
        end
      endcase
    end else begin
      weav_5_8 = 1'b0;
    end
  end

  assign when_Weight_l279_89 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_89) begin
            weav_5_9 = 1'b1;
          end else begin
            weav_5_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_89) begin
            weav_5_9 = 1'b1;
          end else begin
            weav_5_9 = 1'b0;
          end
        end
        default : begin
          weav_5_9 = 1'b0;
        end
      endcase
    end else begin
      weav_5_9 = 1'b0;
    end
  end

  assign when_Weight_l279_90 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_90) begin
            weav_5_10 = 1'b1;
          end else begin
            weav_5_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_90) begin
            weav_5_10 = 1'b1;
          end else begin
            weav_5_10 = 1'b0;
          end
        end
        default : begin
          weav_5_10 = 1'b0;
        end
      endcase
    end else begin
      weav_5_10 = 1'b0;
    end
  end

  assign when_Weight_l279_91 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_91) begin
            weav_5_11 = 1'b1;
          end else begin
            weav_5_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_91) begin
            weav_5_11 = 1'b1;
          end else begin
            weav_5_11 = 1'b0;
          end
        end
        default : begin
          weav_5_11 = 1'b0;
        end
      endcase
    end else begin
      weav_5_11 = 1'b0;
    end
  end

  assign when_Weight_l279_92 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_92) begin
            weav_5_12 = 1'b1;
          end else begin
            weav_5_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_92) begin
            weav_5_12 = 1'b1;
          end else begin
            weav_5_12 = 1'b0;
          end
        end
        default : begin
          weav_5_12 = 1'b0;
        end
      endcase
    end else begin
      weav_5_12 = 1'b0;
    end
  end

  assign when_Weight_l279_93 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_93) begin
            weav_5_13 = 1'b1;
          end else begin
            weav_5_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_93) begin
            weav_5_13 = 1'b1;
          end else begin
            weav_5_13 = 1'b0;
          end
        end
        default : begin
          weav_5_13 = 1'b0;
        end
      endcase
    end else begin
      weav_5_13 = 1'b0;
    end
  end

  assign when_Weight_l279_94 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_94) begin
            weav_5_14 = 1'b1;
          end else begin
            weav_5_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_94) begin
            weav_5_14 = 1'b1;
          end else begin
            weav_5_14 = 1'b0;
          end
        end
        default : begin
          weav_5_14 = 1'b0;
        end
      endcase
    end else begin
      weav_5_14 = 1'b0;
    end
  end

  assign when_Weight_l279_95 = ((copyWeightTimes_count == 4'b0101) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_95) begin
            weav_5_15 = 1'b1;
          end else begin
            weav_5_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_5_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_95) begin
            weav_5_15 = 1'b1;
          end else begin
            weav_5_15 = 1'b0;
          end
        end
        default : begin
          weav_5_15 = 1'b0;
        end
      endcase
    end else begin
      weav_5_15 = 1'b0;
    end
  end

  assign when_Weight_l279_96 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_96) begin
            weav_6_0 = 1'b1;
          end else begin
            weav_6_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_96) begin
            weav_6_0 = 1'b1;
          end else begin
            weav_6_0 = 1'b0;
          end
        end
        default : begin
          weav_6_0 = 1'b0;
        end
      endcase
    end else begin
      weav_6_0 = 1'b0;
    end
  end

  assign when_Weight_l279_97 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_97) begin
            weav_6_1 = 1'b1;
          end else begin
            weav_6_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_97) begin
            weav_6_1 = 1'b1;
          end else begin
            weav_6_1 = 1'b0;
          end
        end
        default : begin
          weav_6_1 = 1'b0;
        end
      endcase
    end else begin
      weav_6_1 = 1'b0;
    end
  end

  assign when_Weight_l279_98 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_98) begin
            weav_6_2 = 1'b1;
          end else begin
            weav_6_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_98) begin
            weav_6_2 = 1'b1;
          end else begin
            weav_6_2 = 1'b0;
          end
        end
        default : begin
          weav_6_2 = 1'b0;
        end
      endcase
    end else begin
      weav_6_2 = 1'b0;
    end
  end

  assign when_Weight_l279_99 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_99) begin
            weav_6_3 = 1'b1;
          end else begin
            weav_6_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_99) begin
            weav_6_3 = 1'b1;
          end else begin
            weav_6_3 = 1'b0;
          end
        end
        default : begin
          weav_6_3 = 1'b0;
        end
      endcase
    end else begin
      weav_6_3 = 1'b0;
    end
  end

  assign when_Weight_l279_100 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_100) begin
            weav_6_4 = 1'b1;
          end else begin
            weav_6_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_100) begin
            weav_6_4 = 1'b1;
          end else begin
            weav_6_4 = 1'b0;
          end
        end
        default : begin
          weav_6_4 = 1'b0;
        end
      endcase
    end else begin
      weav_6_4 = 1'b0;
    end
  end

  assign when_Weight_l279_101 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_101) begin
            weav_6_5 = 1'b1;
          end else begin
            weav_6_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_101) begin
            weav_6_5 = 1'b1;
          end else begin
            weav_6_5 = 1'b0;
          end
        end
        default : begin
          weav_6_5 = 1'b0;
        end
      endcase
    end else begin
      weav_6_5 = 1'b0;
    end
  end

  assign when_Weight_l279_102 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_102) begin
            weav_6_6 = 1'b1;
          end else begin
            weav_6_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_102) begin
            weav_6_6 = 1'b1;
          end else begin
            weav_6_6 = 1'b0;
          end
        end
        default : begin
          weav_6_6 = 1'b0;
        end
      endcase
    end else begin
      weav_6_6 = 1'b0;
    end
  end

  assign when_Weight_l279_103 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_103) begin
            weav_6_7 = 1'b1;
          end else begin
            weav_6_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_103) begin
            weav_6_7 = 1'b1;
          end else begin
            weav_6_7 = 1'b0;
          end
        end
        default : begin
          weav_6_7 = 1'b0;
        end
      endcase
    end else begin
      weav_6_7 = 1'b0;
    end
  end

  assign when_Weight_l279_104 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_104) begin
            weav_6_8 = 1'b1;
          end else begin
            weav_6_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_104) begin
            weav_6_8 = 1'b1;
          end else begin
            weav_6_8 = 1'b0;
          end
        end
        default : begin
          weav_6_8 = 1'b0;
        end
      endcase
    end else begin
      weav_6_8 = 1'b0;
    end
  end

  assign when_Weight_l279_105 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_105) begin
            weav_6_9 = 1'b1;
          end else begin
            weav_6_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_105) begin
            weav_6_9 = 1'b1;
          end else begin
            weav_6_9 = 1'b0;
          end
        end
        default : begin
          weav_6_9 = 1'b0;
        end
      endcase
    end else begin
      weav_6_9 = 1'b0;
    end
  end

  assign when_Weight_l279_106 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_106) begin
            weav_6_10 = 1'b1;
          end else begin
            weav_6_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_106) begin
            weav_6_10 = 1'b1;
          end else begin
            weav_6_10 = 1'b0;
          end
        end
        default : begin
          weav_6_10 = 1'b0;
        end
      endcase
    end else begin
      weav_6_10 = 1'b0;
    end
  end

  assign when_Weight_l279_107 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_107) begin
            weav_6_11 = 1'b1;
          end else begin
            weav_6_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_107) begin
            weav_6_11 = 1'b1;
          end else begin
            weav_6_11 = 1'b0;
          end
        end
        default : begin
          weav_6_11 = 1'b0;
        end
      endcase
    end else begin
      weav_6_11 = 1'b0;
    end
  end

  assign when_Weight_l279_108 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_108) begin
            weav_6_12 = 1'b1;
          end else begin
            weav_6_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_108) begin
            weav_6_12 = 1'b1;
          end else begin
            weav_6_12 = 1'b0;
          end
        end
        default : begin
          weav_6_12 = 1'b0;
        end
      endcase
    end else begin
      weav_6_12 = 1'b0;
    end
  end

  assign when_Weight_l279_109 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_109) begin
            weav_6_13 = 1'b1;
          end else begin
            weav_6_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_109) begin
            weav_6_13 = 1'b1;
          end else begin
            weav_6_13 = 1'b0;
          end
        end
        default : begin
          weav_6_13 = 1'b0;
        end
      endcase
    end else begin
      weav_6_13 = 1'b0;
    end
  end

  assign when_Weight_l279_110 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_110) begin
            weav_6_14 = 1'b1;
          end else begin
            weav_6_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_110) begin
            weav_6_14 = 1'b1;
          end else begin
            weav_6_14 = 1'b0;
          end
        end
        default : begin
          weav_6_14 = 1'b0;
        end
      endcase
    end else begin
      weav_6_14 = 1'b0;
    end
  end

  assign when_Weight_l279_111 = ((copyWeightTimes_count == 4'b0110) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_111) begin
            weav_6_15 = 1'b1;
          end else begin
            weav_6_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_6_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_111) begin
            weav_6_15 = 1'b1;
          end else begin
            weav_6_15 = 1'b0;
          end
        end
        default : begin
          weav_6_15 = 1'b0;
        end
      endcase
    end else begin
      weav_6_15 = 1'b0;
    end
  end

  assign when_Weight_l279_112 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_112) begin
            weav_7_0 = 1'b1;
          end else begin
            weav_7_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_0 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_112) begin
            weav_7_0 = 1'b1;
          end else begin
            weav_7_0 = 1'b0;
          end
        end
        default : begin
          weav_7_0 = 1'b0;
        end
      endcase
    end else begin
      weav_7_0 = 1'b0;
    end
  end

  assign when_Weight_l279_113 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_113) begin
            weav_7_1 = 1'b1;
          end else begin
            weav_7_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_1 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_113) begin
            weav_7_1 = 1'b1;
          end else begin
            weav_7_1 = 1'b0;
          end
        end
        default : begin
          weav_7_1 = 1'b0;
        end
      endcase
    end else begin
      weav_7_1 = 1'b0;
    end
  end

  assign when_Weight_l279_114 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_114) begin
            weav_7_2 = 1'b1;
          end else begin
            weav_7_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_2 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_114) begin
            weav_7_2 = 1'b1;
          end else begin
            weav_7_2 = 1'b0;
          end
        end
        default : begin
          weav_7_2 = 1'b0;
        end
      endcase
    end else begin
      weav_7_2 = 1'b0;
    end
  end

  assign when_Weight_l279_115 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_115) begin
            weav_7_3 = 1'b1;
          end else begin
            weav_7_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_3 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_115) begin
            weav_7_3 = 1'b1;
          end else begin
            weav_7_3 = 1'b0;
          end
        end
        default : begin
          weav_7_3 = 1'b0;
        end
      endcase
    end else begin
      weav_7_3 = 1'b0;
    end
  end

  assign when_Weight_l279_116 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_116) begin
            weav_7_4 = 1'b1;
          end else begin
            weav_7_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_4 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_116) begin
            weav_7_4 = 1'b1;
          end else begin
            weav_7_4 = 1'b0;
          end
        end
        default : begin
          weav_7_4 = 1'b0;
        end
      endcase
    end else begin
      weav_7_4 = 1'b0;
    end
  end

  assign when_Weight_l279_117 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_117) begin
            weav_7_5 = 1'b1;
          end else begin
            weav_7_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_5 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_117) begin
            weav_7_5 = 1'b1;
          end else begin
            weav_7_5 = 1'b0;
          end
        end
        default : begin
          weav_7_5 = 1'b0;
        end
      endcase
    end else begin
      weav_7_5 = 1'b0;
    end
  end

  assign when_Weight_l279_118 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_118) begin
            weav_7_6 = 1'b1;
          end else begin
            weav_7_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_6 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_118) begin
            weav_7_6 = 1'b1;
          end else begin
            weav_7_6 = 1'b0;
          end
        end
        default : begin
          weav_7_6 = 1'b0;
        end
      endcase
    end else begin
      weav_7_6 = 1'b0;
    end
  end

  assign when_Weight_l279_119 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_119) begin
            weav_7_7 = 1'b1;
          end else begin
            weav_7_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_7 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_119) begin
            weav_7_7 = 1'b1;
          end else begin
            weav_7_7 = 1'b0;
          end
        end
        default : begin
          weav_7_7 = 1'b0;
        end
      endcase
    end else begin
      weav_7_7 = 1'b0;
    end
  end

  assign when_Weight_l279_120 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_120) begin
            weav_7_8 = 1'b1;
          end else begin
            weav_7_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_8 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_120) begin
            weav_7_8 = 1'b1;
          end else begin
            weav_7_8 = 1'b0;
          end
        end
        default : begin
          weav_7_8 = 1'b0;
        end
      endcase
    end else begin
      weav_7_8 = 1'b0;
    end
  end

  assign when_Weight_l279_121 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_121) begin
            weav_7_9 = 1'b1;
          end else begin
            weav_7_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_9 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_121) begin
            weav_7_9 = 1'b1;
          end else begin
            weav_7_9 = 1'b0;
          end
        end
        default : begin
          weav_7_9 = 1'b0;
        end
      endcase
    end else begin
      weav_7_9 = 1'b0;
    end
  end

  assign when_Weight_l279_122 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_122) begin
            weav_7_10 = 1'b1;
          end else begin
            weav_7_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_10 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_122) begin
            weav_7_10 = 1'b1;
          end else begin
            weav_7_10 = 1'b0;
          end
        end
        default : begin
          weav_7_10 = 1'b0;
        end
      endcase
    end else begin
      weav_7_10 = 1'b0;
    end
  end

  assign when_Weight_l279_123 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_123) begin
            weav_7_11 = 1'b1;
          end else begin
            weav_7_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_11 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_123) begin
            weav_7_11 = 1'b1;
          end else begin
            weav_7_11 = 1'b0;
          end
        end
        default : begin
          weav_7_11 = 1'b0;
        end
      endcase
    end else begin
      weav_7_11 = 1'b0;
    end
  end

  assign when_Weight_l279_124 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_124) begin
            weav_7_12 = 1'b1;
          end else begin
            weav_7_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_12 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_124) begin
            weav_7_12 = 1'b1;
          end else begin
            weav_7_12 = 1'b0;
          end
        end
        default : begin
          weav_7_12 = 1'b0;
        end
      endcase
    end else begin
      weav_7_12 = 1'b0;
    end
  end

  assign when_Weight_l279_125 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_125) begin
            weav_7_13 = 1'b1;
          end else begin
            weav_7_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_13 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_125) begin
            weav_7_13 = 1'b1;
          end else begin
            weav_7_13 = 1'b0;
          end
        end
        default : begin
          weav_7_13 = 1'b0;
        end
      endcase
    end else begin
      weav_7_13 = 1'b0;
    end
  end

  assign when_Weight_l279_126 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_126) begin
            weav_7_14 = 1'b1;
          end else begin
            weav_7_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_14 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_126) begin
            weav_7_14 = 1'b1;
          end else begin
            weav_7_14 = 1'b0;
          end
        end
        default : begin
          weav_7_14 = 1'b0;
        end
      endcase
    end else begin
      weav_7_14 = 1'b0;
    end
  end

  assign when_Weight_l279_127 = ((copyWeightTimes_count == 4'b0111) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_127) begin
            weav_7_15 = 1'b1;
          end else begin
            weav_7_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_7_15 = 1'b0;
        end
        2'b01 : begin
          if(when_Weight_l306_127) begin
            weav_7_15 = 1'b1;
          end else begin
            weav_7_15 = 1'b0;
          end
        end
        default : begin
          weav_7_15 = 1'b0;
        end
      endcase
    end else begin
      weav_7_15 = 1'b0;
    end
  end

  assign when_Weight_l279_128 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_128) begin
            weav_8_0 = 1'b1;
          end else begin
            weav_8_0 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_0 = 1'b0;
        end
        2'b01 : begin
          weav_8_0 = 1'b0;
        end
        default : begin
          weav_8_0 = 1'b0;
        end
      endcase
    end else begin
      weav_8_0 = 1'b0;
    end
  end

  assign when_Weight_l279_129 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_129) begin
            weav_8_1 = 1'b1;
          end else begin
            weav_8_1 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_1 = 1'b0;
        end
        2'b01 : begin
          weav_8_1 = 1'b0;
        end
        default : begin
          weav_8_1 = 1'b0;
        end
      endcase
    end else begin
      weav_8_1 = 1'b0;
    end
  end

  assign when_Weight_l279_130 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_130) begin
            weav_8_2 = 1'b1;
          end else begin
            weav_8_2 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_2 = 1'b0;
        end
        2'b01 : begin
          weav_8_2 = 1'b0;
        end
        default : begin
          weav_8_2 = 1'b0;
        end
      endcase
    end else begin
      weav_8_2 = 1'b0;
    end
  end

  assign when_Weight_l279_131 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_131) begin
            weav_8_3 = 1'b1;
          end else begin
            weav_8_3 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_3 = 1'b0;
        end
        2'b01 : begin
          weav_8_3 = 1'b0;
        end
        default : begin
          weav_8_3 = 1'b0;
        end
      endcase
    end else begin
      weav_8_3 = 1'b0;
    end
  end

  assign when_Weight_l279_132 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_132) begin
            weav_8_4 = 1'b1;
          end else begin
            weav_8_4 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_4 = 1'b0;
        end
        2'b01 : begin
          weav_8_4 = 1'b0;
        end
        default : begin
          weav_8_4 = 1'b0;
        end
      endcase
    end else begin
      weav_8_4 = 1'b0;
    end
  end

  assign when_Weight_l279_133 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_133) begin
            weav_8_5 = 1'b1;
          end else begin
            weav_8_5 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_5 = 1'b0;
        end
        2'b01 : begin
          weav_8_5 = 1'b0;
        end
        default : begin
          weav_8_5 = 1'b0;
        end
      endcase
    end else begin
      weav_8_5 = 1'b0;
    end
  end

  assign when_Weight_l279_134 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_134) begin
            weav_8_6 = 1'b1;
          end else begin
            weav_8_6 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_6 = 1'b0;
        end
        2'b01 : begin
          weav_8_6 = 1'b0;
        end
        default : begin
          weav_8_6 = 1'b0;
        end
      endcase
    end else begin
      weav_8_6 = 1'b0;
    end
  end

  assign when_Weight_l279_135 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b0111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_135) begin
            weav_8_7 = 1'b1;
          end else begin
            weav_8_7 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_7 = 1'b0;
        end
        2'b01 : begin
          weav_8_7 = 1'b0;
        end
        default : begin
          weav_8_7 = 1'b0;
        end
      endcase
    end else begin
      weav_8_7 = 1'b0;
    end
  end

  assign when_Weight_l279_136 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1000));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_136) begin
            weav_8_8 = 1'b1;
          end else begin
            weav_8_8 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_8 = 1'b0;
        end
        2'b01 : begin
          weav_8_8 = 1'b0;
        end
        default : begin
          weav_8_8 = 1'b0;
        end
      endcase
    end else begin
      weav_8_8 = 1'b0;
    end
  end

  assign when_Weight_l279_137 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1001));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_137) begin
            weav_8_9 = 1'b1;
          end else begin
            weav_8_9 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_9 = 1'b0;
        end
        2'b01 : begin
          weav_8_9 = 1'b0;
        end
        default : begin
          weav_8_9 = 1'b0;
        end
      endcase
    end else begin
      weav_8_9 = 1'b0;
    end
  end

  assign when_Weight_l279_138 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1010));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_138) begin
            weav_8_10 = 1'b1;
          end else begin
            weav_8_10 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_10 = 1'b0;
        end
        2'b01 : begin
          weav_8_10 = 1'b0;
        end
        default : begin
          weav_8_10 = 1'b0;
        end
      endcase
    end else begin
      weav_8_10 = 1'b0;
    end
  end

  assign when_Weight_l279_139 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1011));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_139) begin
            weav_8_11 = 1'b1;
          end else begin
            weav_8_11 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_11 = 1'b0;
        end
        2'b01 : begin
          weav_8_11 = 1'b0;
        end
        default : begin
          weav_8_11 = 1'b0;
        end
      endcase
    end else begin
      weav_8_11 = 1'b0;
    end
  end

  assign when_Weight_l279_140 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1100));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_140) begin
            weav_8_12 = 1'b1;
          end else begin
            weav_8_12 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_12 = 1'b0;
        end
        2'b01 : begin
          weav_8_12 = 1'b0;
        end
        default : begin
          weav_8_12 = 1'b0;
        end
      endcase
    end else begin
      weav_8_12 = 1'b0;
    end
  end

  assign when_Weight_l279_141 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1101));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_141) begin
            weav_8_13 = 1'b1;
          end else begin
            weav_8_13 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_13 = 1'b0;
        end
        2'b01 : begin
          weav_8_13 = 1'b0;
        end
        default : begin
          weav_8_13 = 1'b0;
        end
      endcase
    end else begin
      weav_8_13 = 1'b0;
    end
  end

  assign when_Weight_l279_142 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1110));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_142) begin
            weav_8_14 = 1'b1;
          end else begin
            weav_8_14 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_14 = 1'b0;
        end
        2'b01 : begin
          weav_8_14 = 1'b0;
        end
        default : begin
          weav_8_14 = 1'b0;
        end
      endcase
    end else begin
      weav_8_14 = 1'b0;
    end
  end

  assign when_Weight_l279_143 = ((copyWeightTimes_count == 4'b1000) && (computeChannelOut_count == 4'b1111));
  always @(*) begin
    if(when_Weight_l274) begin
      case(convType)
        2'b00 : begin
          if(when_Weight_l279_143) begin
            weav_8_15 = 1'b1;
          end else begin
            weav_8_15 = 1'b0;
          end
        end
        2'b10 : begin
          weav_8_15 = 1'b0;
        end
        2'b01 : begin
          weav_8_15 = 1'b0;
        end
        default : begin
          weav_8_15 = 1'b0;
        end
      endcase
    end else begin
      weav_8_15 = 1'b0;
    end
  end

  assign when_Weight_l296 = (computeChannelOut_count == 4'b0000);
  assign when_Weight_l296_1 = (computeChannelOut_count == 4'b0001);
  assign when_Weight_l296_2 = (computeChannelOut_count == 4'b0010);
  assign when_Weight_l296_3 = (computeChannelOut_count == 4'b0011);
  assign when_Weight_l296_4 = (computeChannelOut_count == 4'b0100);
  assign when_Weight_l296_5 = (computeChannelOut_count == 4'b0101);
  assign when_Weight_l296_6 = (computeChannelOut_count == 4'b0110);
  assign when_Weight_l296_7 = (computeChannelOut_count == 4'b0111);
  assign when_Weight_l296_8 = (computeChannelOut_count == 4'b1000);
  assign when_Weight_l296_9 = (computeChannelOut_count == 4'b1001);
  assign when_Weight_l296_10 = (computeChannelOut_count == 4'b1010);
  assign when_Weight_l296_11 = (computeChannelOut_count == 4'b1011);
  assign when_Weight_l296_12 = (computeChannelOut_count == 4'b1100);
  assign when_Weight_l296_13 = (computeChannelOut_count == 4'b1101);
  assign when_Weight_l296_14 = (computeChannelOut_count == 4'b1110);
  assign when_Weight_l296_15 = (computeChannelOut_count == 4'b1111);
  assign when_Weight_l306 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_1 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_2 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_3 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_4 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_5 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_6 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_7 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_8 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_9 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_10 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_11 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_12 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_13 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_14 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_15 = ((times_count == 4'b0000) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_16 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_17 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_18 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_19 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_20 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_21 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_22 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_23 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_24 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_25 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_26 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_27 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_28 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_29 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_30 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_31 = ((times_count == 4'b0001) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_32 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_33 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_34 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_35 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_36 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_37 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_38 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_39 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_40 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_41 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_42 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_43 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_44 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_45 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_46 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_47 = ((times_count == 4'b0010) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_48 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_49 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_50 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_51 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_52 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_53 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_54 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_55 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_56 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_57 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_58 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_59 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_60 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_61 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_62 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_63 = ((times_count == 4'b0011) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_64 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_65 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_66 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_67 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_68 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_69 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_70 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_71 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_72 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_73 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_74 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_75 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_76 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_77 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_78 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_79 = ((times_count == 4'b0100) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_80 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_81 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_82 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_83 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_84 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_85 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_86 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_87 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_88 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_89 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_90 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_91 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_92 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_93 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_94 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_95 = ((times_count == 4'b0101) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_96 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_97 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_98 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_99 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_100 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_101 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_102 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_103 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_104 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_105 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_106 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_107 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_108 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_109 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_110 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_111 = ((times_count == 4'b0110) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l306_112 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0000));
  assign when_Weight_l306_113 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0001));
  assign when_Weight_l306_114 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0010));
  assign when_Weight_l306_115 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0011));
  assign when_Weight_l306_116 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0100));
  assign when_Weight_l306_117 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0101));
  assign when_Weight_l306_118 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0110));
  assign when_Weight_l306_119 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b0111));
  assign when_Weight_l306_120 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1000));
  assign when_Weight_l306_121 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1001));
  assign when_Weight_l306_122 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1010));
  assign when_Weight_l306_123 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1011));
  assign when_Weight_l306_124 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1100));
  assign when_Weight_l306_125 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1101));
  assign when_Weight_l306_126 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1110));
  assign when_Weight_l306_127 = ((times_count == 4'b0111) && (computeChannelOut_count == 4'b1111));
  assign when_Weight_l326 = (addr_0_0 == _zz_when_Weight_l326);
  assign when_Weight_l326_1 = (addr_0_1 == _zz_when_Weight_l326_1);
  assign when_Weight_l326_2 = (addr_0_2 == _zz_when_Weight_l326_2);
  assign when_Weight_l326_3 = (addr_0_3 == _zz_when_Weight_l326_3);
  assign when_Weight_l326_4 = (addr_0_4 == _zz_when_Weight_l326_4);
  assign when_Weight_l326_5 = (addr_0_5 == _zz_when_Weight_l326_5);
  assign when_Weight_l326_6 = (addr_0_6 == _zz_when_Weight_l326_6);
  assign when_Weight_l326_7 = (addr_0_7 == _zz_when_Weight_l326_7);
  assign when_Weight_l326_8 = (addr_0_8 == _zz_when_Weight_l326_8);
  assign when_Weight_l326_9 = (addr_0_9 == _zz_when_Weight_l326_9);
  assign when_Weight_l326_10 = (addr_0_10 == _zz_when_Weight_l326_10);
  assign when_Weight_l326_11 = (addr_0_11 == _zz_when_Weight_l326_11);
  assign when_Weight_l326_12 = (addr_0_12 == _zz_when_Weight_l326_12);
  assign when_Weight_l326_13 = (addr_0_13 == _zz_when_Weight_l326_13);
  assign when_Weight_l326_14 = (addr_0_14 == _zz_when_Weight_l326_14);
  assign when_Weight_l326_15 = (addr_0_15 == _zz_when_Weight_l326_15);
  assign when_Weight_l326_16 = (addr_1_0 == _zz_when_Weight_l326_16);
  assign when_Weight_l326_17 = (addr_1_1 == _zz_when_Weight_l326_17);
  assign when_Weight_l326_18 = (addr_1_2 == _zz_when_Weight_l326_18);
  assign when_Weight_l326_19 = (addr_1_3 == _zz_when_Weight_l326_19);
  assign when_Weight_l326_20 = (addr_1_4 == _zz_when_Weight_l326_20);
  assign when_Weight_l326_21 = (addr_1_5 == _zz_when_Weight_l326_21);
  assign when_Weight_l326_22 = (addr_1_6 == _zz_when_Weight_l326_22);
  assign when_Weight_l326_23 = (addr_1_7 == _zz_when_Weight_l326_23);
  assign when_Weight_l326_24 = (addr_1_8 == _zz_when_Weight_l326_24);
  assign when_Weight_l326_25 = (addr_1_9 == _zz_when_Weight_l326_25);
  assign when_Weight_l326_26 = (addr_1_10 == _zz_when_Weight_l326_26);
  assign when_Weight_l326_27 = (addr_1_11 == _zz_when_Weight_l326_27);
  assign when_Weight_l326_28 = (addr_1_12 == _zz_when_Weight_l326_28);
  assign when_Weight_l326_29 = (addr_1_13 == _zz_when_Weight_l326_29);
  assign when_Weight_l326_30 = (addr_1_14 == _zz_when_Weight_l326_30);
  assign when_Weight_l326_31 = (addr_1_15 == _zz_when_Weight_l326_31);
  assign when_Weight_l326_32 = (addr_2_0 == _zz_when_Weight_l326_32);
  assign when_Weight_l326_33 = (addr_2_1 == _zz_when_Weight_l326_33);
  assign when_Weight_l326_34 = (addr_2_2 == _zz_when_Weight_l326_34);
  assign when_Weight_l326_35 = (addr_2_3 == _zz_when_Weight_l326_35);
  assign when_Weight_l326_36 = (addr_2_4 == _zz_when_Weight_l326_36);
  assign when_Weight_l326_37 = (addr_2_5 == _zz_when_Weight_l326_37);
  assign when_Weight_l326_38 = (addr_2_6 == _zz_when_Weight_l326_38);
  assign when_Weight_l326_39 = (addr_2_7 == _zz_when_Weight_l326_39);
  assign when_Weight_l326_40 = (addr_2_8 == _zz_when_Weight_l326_40);
  assign when_Weight_l326_41 = (addr_2_9 == _zz_when_Weight_l326_41);
  assign when_Weight_l326_42 = (addr_2_10 == _zz_when_Weight_l326_42);
  assign when_Weight_l326_43 = (addr_2_11 == _zz_when_Weight_l326_43);
  assign when_Weight_l326_44 = (addr_2_12 == _zz_when_Weight_l326_44);
  assign when_Weight_l326_45 = (addr_2_13 == _zz_when_Weight_l326_45);
  assign when_Weight_l326_46 = (addr_2_14 == _zz_when_Weight_l326_46);
  assign when_Weight_l326_47 = (addr_2_15 == _zz_when_Weight_l326_47);
  assign when_Weight_l326_48 = (addr_3_0 == _zz_when_Weight_l326_48);
  assign when_Weight_l326_49 = (addr_3_1 == _zz_when_Weight_l326_49);
  assign when_Weight_l326_50 = (addr_3_2 == _zz_when_Weight_l326_50);
  assign when_Weight_l326_51 = (addr_3_3 == _zz_when_Weight_l326_51);
  assign when_Weight_l326_52 = (addr_3_4 == _zz_when_Weight_l326_52);
  assign when_Weight_l326_53 = (addr_3_5 == _zz_when_Weight_l326_53);
  assign when_Weight_l326_54 = (addr_3_6 == _zz_when_Weight_l326_54);
  assign when_Weight_l326_55 = (addr_3_7 == _zz_when_Weight_l326_55);
  assign when_Weight_l326_56 = (addr_3_8 == _zz_when_Weight_l326_56);
  assign when_Weight_l326_57 = (addr_3_9 == _zz_when_Weight_l326_57);
  assign when_Weight_l326_58 = (addr_3_10 == _zz_when_Weight_l326_58);
  assign when_Weight_l326_59 = (addr_3_11 == _zz_when_Weight_l326_59);
  assign when_Weight_l326_60 = (addr_3_12 == _zz_when_Weight_l326_60);
  assign when_Weight_l326_61 = (addr_3_13 == _zz_when_Weight_l326_61);
  assign when_Weight_l326_62 = (addr_3_14 == _zz_when_Weight_l326_62);
  assign when_Weight_l326_63 = (addr_3_15 == _zz_when_Weight_l326_63);
  assign when_Weight_l326_64 = (addr_4_0 == _zz_when_Weight_l326_64);
  assign when_Weight_l326_65 = (addr_4_1 == _zz_when_Weight_l326_65);
  assign when_Weight_l326_66 = (addr_4_2 == _zz_when_Weight_l326_66);
  assign when_Weight_l326_67 = (addr_4_3 == _zz_when_Weight_l326_67);
  assign when_Weight_l326_68 = (addr_4_4 == _zz_when_Weight_l326_68);
  assign when_Weight_l326_69 = (addr_4_5 == _zz_when_Weight_l326_69);
  assign when_Weight_l326_70 = (addr_4_6 == _zz_when_Weight_l326_70);
  assign when_Weight_l326_71 = (addr_4_7 == _zz_when_Weight_l326_71);
  assign when_Weight_l326_72 = (addr_4_8 == _zz_when_Weight_l326_72);
  assign when_Weight_l326_73 = (addr_4_9 == _zz_when_Weight_l326_73);
  assign when_Weight_l326_74 = (addr_4_10 == _zz_when_Weight_l326_74);
  assign when_Weight_l326_75 = (addr_4_11 == _zz_when_Weight_l326_75);
  assign when_Weight_l326_76 = (addr_4_12 == _zz_when_Weight_l326_76);
  assign when_Weight_l326_77 = (addr_4_13 == _zz_when_Weight_l326_77);
  assign when_Weight_l326_78 = (addr_4_14 == _zz_when_Weight_l326_78);
  assign when_Weight_l326_79 = (addr_4_15 == _zz_when_Weight_l326_79);
  assign when_Weight_l326_80 = (addr_5_0 == _zz_when_Weight_l326_80);
  assign when_Weight_l326_81 = (addr_5_1 == _zz_when_Weight_l326_81);
  assign when_Weight_l326_82 = (addr_5_2 == _zz_when_Weight_l326_82);
  assign when_Weight_l326_83 = (addr_5_3 == _zz_when_Weight_l326_83);
  assign when_Weight_l326_84 = (addr_5_4 == _zz_when_Weight_l326_84);
  assign when_Weight_l326_85 = (addr_5_5 == _zz_when_Weight_l326_85);
  assign when_Weight_l326_86 = (addr_5_6 == _zz_when_Weight_l326_86);
  assign when_Weight_l326_87 = (addr_5_7 == _zz_when_Weight_l326_87);
  assign when_Weight_l326_88 = (addr_5_8 == _zz_when_Weight_l326_88);
  assign when_Weight_l326_89 = (addr_5_9 == _zz_when_Weight_l326_89);
  assign when_Weight_l326_90 = (addr_5_10 == _zz_when_Weight_l326_90);
  assign when_Weight_l326_91 = (addr_5_11 == _zz_when_Weight_l326_91);
  assign when_Weight_l326_92 = (addr_5_12 == _zz_when_Weight_l326_92);
  assign when_Weight_l326_93 = (addr_5_13 == _zz_when_Weight_l326_93);
  assign when_Weight_l326_94 = (addr_5_14 == _zz_when_Weight_l326_94);
  assign when_Weight_l326_95 = (addr_5_15 == _zz_when_Weight_l326_95);
  assign when_Weight_l326_96 = (addr_6_0 == _zz_when_Weight_l326_96);
  assign when_Weight_l326_97 = (addr_6_1 == _zz_when_Weight_l326_97);
  assign when_Weight_l326_98 = (addr_6_2 == _zz_when_Weight_l326_98);
  assign when_Weight_l326_99 = (addr_6_3 == _zz_when_Weight_l326_99);
  assign when_Weight_l326_100 = (addr_6_4 == _zz_when_Weight_l326_100);
  assign when_Weight_l326_101 = (addr_6_5 == _zz_when_Weight_l326_101);
  assign when_Weight_l326_102 = (addr_6_6 == _zz_when_Weight_l326_102);
  assign when_Weight_l326_103 = (addr_6_7 == _zz_when_Weight_l326_103);
  assign when_Weight_l326_104 = (addr_6_8 == _zz_when_Weight_l326_104);
  assign when_Weight_l326_105 = (addr_6_9 == _zz_when_Weight_l326_105);
  assign when_Weight_l326_106 = (addr_6_10 == _zz_when_Weight_l326_106);
  assign when_Weight_l326_107 = (addr_6_11 == _zz_when_Weight_l326_107);
  assign when_Weight_l326_108 = (addr_6_12 == _zz_when_Weight_l326_108);
  assign when_Weight_l326_109 = (addr_6_13 == _zz_when_Weight_l326_109);
  assign when_Weight_l326_110 = (addr_6_14 == _zz_when_Weight_l326_110);
  assign when_Weight_l326_111 = (addr_6_15 == _zz_when_Weight_l326_111);
  assign when_Weight_l326_112 = (addr_7_0 == _zz_when_Weight_l326_112);
  assign when_Weight_l326_113 = (addr_7_1 == _zz_when_Weight_l326_113);
  assign when_Weight_l326_114 = (addr_7_2 == _zz_when_Weight_l326_114);
  assign when_Weight_l326_115 = (addr_7_3 == _zz_when_Weight_l326_115);
  assign when_Weight_l326_116 = (addr_7_4 == _zz_when_Weight_l326_116);
  assign when_Weight_l326_117 = (addr_7_5 == _zz_when_Weight_l326_117);
  assign when_Weight_l326_118 = (addr_7_6 == _zz_when_Weight_l326_118);
  assign when_Weight_l326_119 = (addr_7_7 == _zz_when_Weight_l326_119);
  assign when_Weight_l326_120 = (addr_7_8 == _zz_when_Weight_l326_120);
  assign when_Weight_l326_121 = (addr_7_9 == _zz_when_Weight_l326_121);
  assign when_Weight_l326_122 = (addr_7_10 == _zz_when_Weight_l326_122);
  assign when_Weight_l326_123 = (addr_7_11 == _zz_when_Weight_l326_123);
  assign when_Weight_l326_124 = (addr_7_12 == _zz_when_Weight_l326_124);
  assign when_Weight_l326_125 = (addr_7_13 == _zz_when_Weight_l326_125);
  assign when_Weight_l326_126 = (addr_7_14 == _zz_when_Weight_l326_126);
  assign when_Weight_l326_127 = (addr_7_15 == _zz_when_Weight_l326_127);
  assign when_Weight_l326_128 = (addr_8_0 == _zz_when_Weight_l326_128);
  assign when_Weight_l326_129 = (addr_8_1 == _zz_when_Weight_l326_129);
  assign when_Weight_l326_130 = (addr_8_2 == _zz_when_Weight_l326_130);
  assign when_Weight_l326_131 = (addr_8_3 == _zz_when_Weight_l326_131);
  assign when_Weight_l326_132 = (addr_8_4 == _zz_when_Weight_l326_132);
  assign when_Weight_l326_133 = (addr_8_5 == _zz_when_Weight_l326_133);
  assign when_Weight_l326_134 = (addr_8_6 == _zz_when_Weight_l326_134);
  assign when_Weight_l326_135 = (addr_8_7 == _zz_when_Weight_l326_135);
  assign when_Weight_l326_136 = (addr_8_8 == _zz_when_Weight_l326_136);
  assign when_Weight_l326_137 = (addr_8_9 == _zz_when_Weight_l326_137);
  assign when_Weight_l326_138 = (addr_8_10 == _zz_when_Weight_l326_138);
  assign when_Weight_l326_139 = (addr_8_11 == _zz_when_Weight_l326_139);
  assign when_Weight_l326_140 = (addr_8_12 == _zz_when_Weight_l326_140);
  assign when_Weight_l326_141 = (addr_8_13 == _zz_when_Weight_l326_141);
  assign when_Weight_l326_142 = (addr_8_14 == _zz_when_Weight_l326_142);
  assign when_Weight_l326_143 = (addr_8_15 == _zz_when_Weight_l326_143);
  assign weightRead_0_data = {{{{{{_zz_weightRead_0_data,weightData_0_5},weightData_0_4},weightData_0_3},weightData_0_2},weightData_0_1},weightData_0_0};
  assign weightRead_1_data = {{{{{{_zz_weightRead_1_data,weightData_1_5},weightData_1_4},weightData_1_3},weightData_1_2},weightData_1_1},weightData_1_0};
  assign weightRead_2_data = {{{{{{_zz_weightRead_2_data,weightData_2_5},weightData_2_4},weightData_2_3},weightData_2_2},weightData_2_1},weightData_2_0};
  assign weightRead_3_data = {{{{{{_zz_weightRead_3_data,weightData_3_5},weightData_3_4},weightData_3_3},weightData_3_2},weightData_3_1},weightData_3_0};
  assign weightRead_4_data = {{{{{{_zz_weightRead_4_data,weightData_4_5},weightData_4_4},weightData_4_3},weightData_4_2},weightData_4_1},weightData_4_0};
  assign weightRead_5_data = {{{{{{_zz_weightRead_5_data,weightData_5_5},weightData_5_4},weightData_5_3},weightData_5_2},weightData_5_1},weightData_5_0};
  assign weightRead_6_data = {{{{{{_zz_weightRead_6_data,weightData_6_5},weightData_6_4},weightData_6_3},weightData_6_2},weightData_6_1},weightData_6_0};
  assign weightRead_7_data = {{{{{{_zz_weightRead_7_data,weightData_7_5},weightData_7_4},weightData_7_3},weightData_7_2},weightData_7_1},weightData_7_0};
  assign weightRead_8_data = {{{{{{_zz_weightRead_8_data,weightData_8_5},weightData_8_4},weightData_8_3},weightData_8_2},weightData_8_1},weightData_8_0};
  assign weightRam_0_0_wea = weav_0_0;
  assign weightRam_0_0_addrb = weightRead_0_addr;
  assign weightData_0_0 = weightRam_0_0_doutb;
  assign weightRam_0_0_addra = _zz_addra[8:0];
  assign weightRam_0_0_dina = sData_payload;
  assign weightRam_0_1_wea = weav_0_1;
  assign weightRam_0_1_addrb = weightRead_0_addr;
  assign weightData_0_1 = weightRam_0_1_doutb;
  assign weightRam_0_1_addra = _zz_addra_1[8:0];
  assign weightRam_0_1_dina = sData_payload;
  assign weightRam_0_2_wea = weav_0_2;
  assign weightRam_0_2_addrb = weightRead_0_addr;
  assign weightData_0_2 = weightRam_0_2_doutb;
  assign weightRam_0_2_addra = _zz_addra_2[8:0];
  assign weightRam_0_2_dina = sData_payload;
  assign weightRam_0_3_wea = weav_0_3;
  assign weightRam_0_3_addrb = weightRead_0_addr;
  assign weightData_0_3 = weightRam_0_3_doutb;
  assign weightRam_0_3_addra = _zz_addra_3[8:0];
  assign weightRam_0_3_dina = sData_payload;
  assign weightRam_0_4_wea = weav_0_4;
  assign weightRam_0_4_addrb = weightRead_0_addr;
  assign weightData_0_4 = weightRam_0_4_doutb;
  assign weightRam_0_4_addra = _zz_addra_4[8:0];
  assign weightRam_0_4_dina = sData_payload;
  assign weightRam_0_5_wea = weav_0_5;
  assign weightRam_0_5_addrb = weightRead_0_addr;
  assign weightData_0_5 = weightRam_0_5_doutb;
  assign weightRam_0_5_addra = _zz_addra_5[8:0];
  assign weightRam_0_5_dina = sData_payload;
  assign weightRam_0_6_wea = weav_0_6;
  assign weightRam_0_6_addrb = weightRead_0_addr;
  assign weightData_0_6 = weightRam_0_6_doutb;
  assign weightRam_0_6_addra = _zz_addra_6[8:0];
  assign weightRam_0_6_dina = sData_payload;
  assign weightRam_0_7_wea = weav_0_7;
  assign weightRam_0_7_addrb = weightRead_0_addr;
  assign weightData_0_7 = weightRam_0_7_doutb;
  assign weightRam_0_7_addra = _zz_addra_7[8:0];
  assign weightRam_0_7_dina = sData_payload;
  assign weightRam_0_8_wea = weav_0_8;
  assign weightRam_0_8_addrb = weightRead_0_addr;
  assign weightData_0_8 = weightRam_0_8_doutb;
  assign weightRam_0_8_addra = _zz_addra_8[8:0];
  assign weightRam_0_8_dina = sData_payload;
  assign weightRam_0_9_wea = weav_0_9;
  assign weightRam_0_9_addrb = weightRead_0_addr;
  assign weightData_0_9 = weightRam_0_9_doutb;
  assign weightRam_0_9_addra = _zz_addra_9[8:0];
  assign weightRam_0_9_dina = sData_payload;
  assign weightRam_0_10_wea = weav_0_10;
  assign weightRam_0_10_addrb = weightRead_0_addr;
  assign weightData_0_10 = weightRam_0_10_doutb;
  assign weightRam_0_10_addra = _zz_addra_10[8:0];
  assign weightRam_0_10_dina = sData_payload;
  assign weightRam_0_11_wea = weav_0_11;
  assign weightRam_0_11_addrb = weightRead_0_addr;
  assign weightData_0_11 = weightRam_0_11_doutb;
  assign weightRam_0_11_addra = _zz_addra_11[8:0];
  assign weightRam_0_11_dina = sData_payload;
  assign weightRam_0_12_wea = weav_0_12;
  assign weightRam_0_12_addrb = weightRead_0_addr;
  assign weightData_0_12 = weightRam_0_12_doutb;
  assign weightRam_0_12_addra = _zz_addra_12[8:0];
  assign weightRam_0_12_dina = sData_payload;
  assign weightRam_0_13_wea = weav_0_13;
  assign weightRam_0_13_addrb = weightRead_0_addr;
  assign weightData_0_13 = weightRam_0_13_doutb;
  assign weightRam_0_13_addra = _zz_addra_13[8:0];
  assign weightRam_0_13_dina = sData_payload;
  assign weightRam_0_14_wea = weav_0_14;
  assign weightRam_0_14_addrb = weightRead_0_addr;
  assign weightData_0_14 = weightRam_0_14_doutb;
  assign weightRam_0_14_addra = _zz_addra_14[8:0];
  assign weightRam_0_14_dina = sData_payload;
  assign weightRam_0_15_wea = weav_0_15;
  assign weightRam_0_15_addrb = weightRead_0_addr;
  assign weightData_0_15 = weightRam_0_15_doutb;
  assign weightRam_0_15_addra = _zz_addra_15[8:0];
  assign weightRam_0_15_dina = sData_payload;
  assign weightRam_1_0_wea = weav_1_0;
  assign weightRam_1_0_addrb = weightRead_1_addr;
  assign weightData_1_0 = weightRam_1_0_doutb;
  assign weightRam_1_0_addra = _zz_addra_16[8:0];
  assign weightRam_1_0_dina = sData_payload;
  assign weightRam_1_1_wea = weav_1_1;
  assign weightRam_1_1_addrb = weightRead_1_addr;
  assign weightData_1_1 = weightRam_1_1_doutb;
  assign weightRam_1_1_addra = _zz_addra_17[8:0];
  assign weightRam_1_1_dina = sData_payload;
  assign weightRam_1_2_wea = weav_1_2;
  assign weightRam_1_2_addrb = weightRead_1_addr;
  assign weightData_1_2 = weightRam_1_2_doutb;
  assign weightRam_1_2_addra = _zz_addra_18[8:0];
  assign weightRam_1_2_dina = sData_payload;
  assign weightRam_1_3_wea = weav_1_3;
  assign weightRam_1_3_addrb = weightRead_1_addr;
  assign weightData_1_3 = weightRam_1_3_doutb;
  assign weightRam_1_3_addra = _zz_addra_19[8:0];
  assign weightRam_1_3_dina = sData_payload;
  assign weightRam_1_4_wea = weav_1_4;
  assign weightRam_1_4_addrb = weightRead_1_addr;
  assign weightData_1_4 = weightRam_1_4_doutb;
  assign weightRam_1_4_addra = _zz_addra_20[8:0];
  assign weightRam_1_4_dina = sData_payload;
  assign weightRam_1_5_wea = weav_1_5;
  assign weightRam_1_5_addrb = weightRead_1_addr;
  assign weightData_1_5 = weightRam_1_5_doutb;
  assign weightRam_1_5_addra = _zz_addra_21[8:0];
  assign weightRam_1_5_dina = sData_payload;
  assign weightRam_1_6_wea = weav_1_6;
  assign weightRam_1_6_addrb = weightRead_1_addr;
  assign weightData_1_6 = weightRam_1_6_doutb;
  assign weightRam_1_6_addra = _zz_addra_22[8:0];
  assign weightRam_1_6_dina = sData_payload;
  assign weightRam_1_7_wea = weav_1_7;
  assign weightRam_1_7_addrb = weightRead_1_addr;
  assign weightData_1_7 = weightRam_1_7_doutb;
  assign weightRam_1_7_addra = _zz_addra_23[8:0];
  assign weightRam_1_7_dina = sData_payload;
  assign weightRam_1_8_wea = weav_1_8;
  assign weightRam_1_8_addrb = weightRead_1_addr;
  assign weightData_1_8 = weightRam_1_8_doutb;
  assign weightRam_1_8_addra = _zz_addra_24[8:0];
  assign weightRam_1_8_dina = sData_payload;
  assign weightRam_1_9_wea = weav_1_9;
  assign weightRam_1_9_addrb = weightRead_1_addr;
  assign weightData_1_9 = weightRam_1_9_doutb;
  assign weightRam_1_9_addra = _zz_addra_25[8:0];
  assign weightRam_1_9_dina = sData_payload;
  assign weightRam_1_10_wea = weav_1_10;
  assign weightRam_1_10_addrb = weightRead_1_addr;
  assign weightData_1_10 = weightRam_1_10_doutb;
  assign weightRam_1_10_addra = _zz_addra_26[8:0];
  assign weightRam_1_10_dina = sData_payload;
  assign weightRam_1_11_wea = weav_1_11;
  assign weightRam_1_11_addrb = weightRead_1_addr;
  assign weightData_1_11 = weightRam_1_11_doutb;
  assign weightRam_1_11_addra = _zz_addra_27[8:0];
  assign weightRam_1_11_dina = sData_payload;
  assign weightRam_1_12_wea = weav_1_12;
  assign weightRam_1_12_addrb = weightRead_1_addr;
  assign weightData_1_12 = weightRam_1_12_doutb;
  assign weightRam_1_12_addra = _zz_addra_28[8:0];
  assign weightRam_1_12_dina = sData_payload;
  assign weightRam_1_13_wea = weav_1_13;
  assign weightRam_1_13_addrb = weightRead_1_addr;
  assign weightData_1_13 = weightRam_1_13_doutb;
  assign weightRam_1_13_addra = _zz_addra_29[8:0];
  assign weightRam_1_13_dina = sData_payload;
  assign weightRam_1_14_wea = weav_1_14;
  assign weightRam_1_14_addrb = weightRead_1_addr;
  assign weightData_1_14 = weightRam_1_14_doutb;
  assign weightRam_1_14_addra = _zz_addra_30[8:0];
  assign weightRam_1_14_dina = sData_payload;
  assign weightRam_1_15_wea = weav_1_15;
  assign weightRam_1_15_addrb = weightRead_1_addr;
  assign weightData_1_15 = weightRam_1_15_doutb;
  assign weightRam_1_15_addra = _zz_addra_31[8:0];
  assign weightRam_1_15_dina = sData_payload;
  assign weightRam_2_0_wea = weav_2_0;
  assign weightRam_2_0_addrb = weightRead_2_addr;
  assign weightData_2_0 = weightRam_2_0_doutb;
  assign weightRam_2_0_addra = _zz_addra_32[8:0];
  assign weightRam_2_0_dina = sData_payload;
  assign weightRam_2_1_wea = weav_2_1;
  assign weightRam_2_1_addrb = weightRead_2_addr;
  assign weightData_2_1 = weightRam_2_1_doutb;
  assign weightRam_2_1_addra = _zz_addra_33[8:0];
  assign weightRam_2_1_dina = sData_payload;
  assign weightRam_2_2_wea = weav_2_2;
  assign weightRam_2_2_addrb = weightRead_2_addr;
  assign weightData_2_2 = weightRam_2_2_doutb;
  assign weightRam_2_2_addra = _zz_addra_34[8:0];
  assign weightRam_2_2_dina = sData_payload;
  assign weightRam_2_3_wea = weav_2_3;
  assign weightRam_2_3_addrb = weightRead_2_addr;
  assign weightData_2_3 = weightRam_2_3_doutb;
  assign weightRam_2_3_addra = _zz_addra_35[8:0];
  assign weightRam_2_3_dina = sData_payload;
  assign weightRam_2_4_wea = weav_2_4;
  assign weightRam_2_4_addrb = weightRead_2_addr;
  assign weightData_2_4 = weightRam_2_4_doutb;
  assign weightRam_2_4_addra = _zz_addra_36[8:0];
  assign weightRam_2_4_dina = sData_payload;
  assign weightRam_2_5_wea = weav_2_5;
  assign weightRam_2_5_addrb = weightRead_2_addr;
  assign weightData_2_5 = weightRam_2_5_doutb;
  assign weightRam_2_5_addra = _zz_addra_37[8:0];
  assign weightRam_2_5_dina = sData_payload;
  assign weightRam_2_6_wea = weav_2_6;
  assign weightRam_2_6_addrb = weightRead_2_addr;
  assign weightData_2_6 = weightRam_2_6_doutb;
  assign weightRam_2_6_addra = _zz_addra_38[8:0];
  assign weightRam_2_6_dina = sData_payload;
  assign weightRam_2_7_wea = weav_2_7;
  assign weightRam_2_7_addrb = weightRead_2_addr;
  assign weightData_2_7 = weightRam_2_7_doutb;
  assign weightRam_2_7_addra = _zz_addra_39[8:0];
  assign weightRam_2_7_dina = sData_payload;
  assign weightRam_2_8_wea = weav_2_8;
  assign weightRam_2_8_addrb = weightRead_2_addr;
  assign weightData_2_8 = weightRam_2_8_doutb;
  assign weightRam_2_8_addra = _zz_addra_40[8:0];
  assign weightRam_2_8_dina = sData_payload;
  assign weightRam_2_9_wea = weav_2_9;
  assign weightRam_2_9_addrb = weightRead_2_addr;
  assign weightData_2_9 = weightRam_2_9_doutb;
  assign weightRam_2_9_addra = _zz_addra_41[8:0];
  assign weightRam_2_9_dina = sData_payload;
  assign weightRam_2_10_wea = weav_2_10;
  assign weightRam_2_10_addrb = weightRead_2_addr;
  assign weightData_2_10 = weightRam_2_10_doutb;
  assign weightRam_2_10_addra = _zz_addra_42[8:0];
  assign weightRam_2_10_dina = sData_payload;
  assign weightRam_2_11_wea = weav_2_11;
  assign weightRam_2_11_addrb = weightRead_2_addr;
  assign weightData_2_11 = weightRam_2_11_doutb;
  assign weightRam_2_11_addra = _zz_addra_43[8:0];
  assign weightRam_2_11_dina = sData_payload;
  assign weightRam_2_12_wea = weav_2_12;
  assign weightRam_2_12_addrb = weightRead_2_addr;
  assign weightData_2_12 = weightRam_2_12_doutb;
  assign weightRam_2_12_addra = _zz_addra_44[8:0];
  assign weightRam_2_12_dina = sData_payload;
  assign weightRam_2_13_wea = weav_2_13;
  assign weightRam_2_13_addrb = weightRead_2_addr;
  assign weightData_2_13 = weightRam_2_13_doutb;
  assign weightRam_2_13_addra = _zz_addra_45[8:0];
  assign weightRam_2_13_dina = sData_payload;
  assign weightRam_2_14_wea = weav_2_14;
  assign weightRam_2_14_addrb = weightRead_2_addr;
  assign weightData_2_14 = weightRam_2_14_doutb;
  assign weightRam_2_14_addra = _zz_addra_46[8:0];
  assign weightRam_2_14_dina = sData_payload;
  assign weightRam_2_15_wea = weav_2_15;
  assign weightRam_2_15_addrb = weightRead_2_addr;
  assign weightData_2_15 = weightRam_2_15_doutb;
  assign weightRam_2_15_addra = _zz_addra_47[8:0];
  assign weightRam_2_15_dina = sData_payload;
  assign weightRam_3_0_wea = weav_3_0;
  assign weightRam_3_0_addrb = weightRead_3_addr;
  assign weightData_3_0 = weightRam_3_0_doutb;
  assign weightRam_3_0_addra = _zz_addra_48[8:0];
  assign weightRam_3_0_dina = sData_payload;
  assign weightRam_3_1_wea = weav_3_1;
  assign weightRam_3_1_addrb = weightRead_3_addr;
  assign weightData_3_1 = weightRam_3_1_doutb;
  assign weightRam_3_1_addra = _zz_addra_49[8:0];
  assign weightRam_3_1_dina = sData_payload;
  assign weightRam_3_2_wea = weav_3_2;
  assign weightRam_3_2_addrb = weightRead_3_addr;
  assign weightData_3_2 = weightRam_3_2_doutb;
  assign weightRam_3_2_addra = _zz_addra_50[8:0];
  assign weightRam_3_2_dina = sData_payload;
  assign weightRam_3_3_wea = weav_3_3;
  assign weightRam_3_3_addrb = weightRead_3_addr;
  assign weightData_3_3 = weightRam_3_3_doutb;
  assign weightRam_3_3_addra = _zz_addra_51[8:0];
  assign weightRam_3_3_dina = sData_payload;
  assign weightRam_3_4_wea = weav_3_4;
  assign weightRam_3_4_addrb = weightRead_3_addr;
  assign weightData_3_4 = weightRam_3_4_doutb;
  assign weightRam_3_4_addra = _zz_addra_52[8:0];
  assign weightRam_3_4_dina = sData_payload;
  assign weightRam_3_5_wea = weav_3_5;
  assign weightRam_3_5_addrb = weightRead_3_addr;
  assign weightData_3_5 = weightRam_3_5_doutb;
  assign weightRam_3_5_addra = _zz_addra_53[8:0];
  assign weightRam_3_5_dina = sData_payload;
  assign weightRam_3_6_wea = weav_3_6;
  assign weightRam_3_6_addrb = weightRead_3_addr;
  assign weightData_3_6 = weightRam_3_6_doutb;
  assign weightRam_3_6_addra = _zz_addra_54[8:0];
  assign weightRam_3_6_dina = sData_payload;
  assign weightRam_3_7_wea = weav_3_7;
  assign weightRam_3_7_addrb = weightRead_3_addr;
  assign weightData_3_7 = weightRam_3_7_doutb;
  assign weightRam_3_7_addra = _zz_addra_55[8:0];
  assign weightRam_3_7_dina = sData_payload;
  assign weightRam_3_8_wea = weav_3_8;
  assign weightRam_3_8_addrb = weightRead_3_addr;
  assign weightData_3_8 = weightRam_3_8_doutb;
  assign weightRam_3_8_addra = _zz_addra_56[8:0];
  assign weightRam_3_8_dina = sData_payload;
  assign weightRam_3_9_wea = weav_3_9;
  assign weightRam_3_9_addrb = weightRead_3_addr;
  assign weightData_3_9 = weightRam_3_9_doutb;
  assign weightRam_3_9_addra = _zz_addra_57[8:0];
  assign weightRam_3_9_dina = sData_payload;
  assign weightRam_3_10_wea = weav_3_10;
  assign weightRam_3_10_addrb = weightRead_3_addr;
  assign weightData_3_10 = weightRam_3_10_doutb;
  assign weightRam_3_10_addra = _zz_addra_58[8:0];
  assign weightRam_3_10_dina = sData_payload;
  assign weightRam_3_11_wea = weav_3_11;
  assign weightRam_3_11_addrb = weightRead_3_addr;
  assign weightData_3_11 = weightRam_3_11_doutb;
  assign weightRam_3_11_addra = _zz_addra_59[8:0];
  assign weightRam_3_11_dina = sData_payload;
  assign weightRam_3_12_wea = weav_3_12;
  assign weightRam_3_12_addrb = weightRead_3_addr;
  assign weightData_3_12 = weightRam_3_12_doutb;
  assign weightRam_3_12_addra = _zz_addra_60[8:0];
  assign weightRam_3_12_dina = sData_payload;
  assign weightRam_3_13_wea = weav_3_13;
  assign weightRam_3_13_addrb = weightRead_3_addr;
  assign weightData_3_13 = weightRam_3_13_doutb;
  assign weightRam_3_13_addra = _zz_addra_61[8:0];
  assign weightRam_3_13_dina = sData_payload;
  assign weightRam_3_14_wea = weav_3_14;
  assign weightRam_3_14_addrb = weightRead_3_addr;
  assign weightData_3_14 = weightRam_3_14_doutb;
  assign weightRam_3_14_addra = _zz_addra_62[8:0];
  assign weightRam_3_14_dina = sData_payload;
  assign weightRam_3_15_wea = weav_3_15;
  assign weightRam_3_15_addrb = weightRead_3_addr;
  assign weightData_3_15 = weightRam_3_15_doutb;
  assign weightRam_3_15_addra = _zz_addra_63[8:0];
  assign weightRam_3_15_dina = sData_payload;
  assign weightRam_4_0_wea = weav_4_0;
  assign weightRam_4_0_addrb = weightRead_4_addr;
  assign weightData_4_0 = weightRam_4_0_doutb;
  assign weightRam_4_0_addra = _zz_addra_64[8:0];
  assign weightRam_4_0_dina = sData_payload;
  assign weightRam_4_1_wea = weav_4_1;
  assign weightRam_4_1_addrb = weightRead_4_addr;
  assign weightData_4_1 = weightRam_4_1_doutb;
  assign weightRam_4_1_addra = _zz_addra_65[8:0];
  assign weightRam_4_1_dina = sData_payload;
  assign weightRam_4_2_wea = weav_4_2;
  assign weightRam_4_2_addrb = weightRead_4_addr;
  assign weightData_4_2 = weightRam_4_2_doutb;
  assign weightRam_4_2_addra = _zz_addra_66[8:0];
  assign weightRam_4_2_dina = sData_payload;
  assign weightRam_4_3_wea = weav_4_3;
  assign weightRam_4_3_addrb = weightRead_4_addr;
  assign weightData_4_3 = weightRam_4_3_doutb;
  assign weightRam_4_3_addra = _zz_addra_67[8:0];
  assign weightRam_4_3_dina = sData_payload;
  assign weightRam_4_4_wea = weav_4_4;
  assign weightRam_4_4_addrb = weightRead_4_addr;
  assign weightData_4_4 = weightRam_4_4_doutb;
  assign weightRam_4_4_addra = _zz_addra_68[8:0];
  assign weightRam_4_4_dina = sData_payload;
  assign weightRam_4_5_wea = weav_4_5;
  assign weightRam_4_5_addrb = weightRead_4_addr;
  assign weightData_4_5 = weightRam_4_5_doutb;
  assign weightRam_4_5_addra = _zz_addra_69[8:0];
  assign weightRam_4_5_dina = sData_payload;
  assign weightRam_4_6_wea = weav_4_6;
  assign weightRam_4_6_addrb = weightRead_4_addr;
  assign weightData_4_6 = weightRam_4_6_doutb;
  assign weightRam_4_6_addra = _zz_addra_70[8:0];
  assign weightRam_4_6_dina = sData_payload;
  assign weightRam_4_7_wea = weav_4_7;
  assign weightRam_4_7_addrb = weightRead_4_addr;
  assign weightData_4_7 = weightRam_4_7_doutb;
  assign weightRam_4_7_addra = _zz_addra_71[8:0];
  assign weightRam_4_7_dina = sData_payload;
  assign weightRam_4_8_wea = weav_4_8;
  assign weightRam_4_8_addrb = weightRead_4_addr;
  assign weightData_4_8 = weightRam_4_8_doutb;
  assign weightRam_4_8_addra = _zz_addra_72[8:0];
  assign weightRam_4_8_dina = sData_payload;
  assign weightRam_4_9_wea = weav_4_9;
  assign weightRam_4_9_addrb = weightRead_4_addr;
  assign weightData_4_9 = weightRam_4_9_doutb;
  assign weightRam_4_9_addra = _zz_addra_73[8:0];
  assign weightRam_4_9_dina = sData_payload;
  assign weightRam_4_10_wea = weav_4_10;
  assign weightRam_4_10_addrb = weightRead_4_addr;
  assign weightData_4_10 = weightRam_4_10_doutb;
  assign weightRam_4_10_addra = _zz_addra_74[8:0];
  assign weightRam_4_10_dina = sData_payload;
  assign weightRam_4_11_wea = weav_4_11;
  assign weightRam_4_11_addrb = weightRead_4_addr;
  assign weightData_4_11 = weightRam_4_11_doutb;
  assign weightRam_4_11_addra = _zz_addra_75[8:0];
  assign weightRam_4_11_dina = sData_payload;
  assign weightRam_4_12_wea = weav_4_12;
  assign weightRam_4_12_addrb = weightRead_4_addr;
  assign weightData_4_12 = weightRam_4_12_doutb;
  assign weightRam_4_12_addra = _zz_addra_76[8:0];
  assign weightRam_4_12_dina = sData_payload;
  assign weightRam_4_13_wea = weav_4_13;
  assign weightRam_4_13_addrb = weightRead_4_addr;
  assign weightData_4_13 = weightRam_4_13_doutb;
  assign weightRam_4_13_addra = _zz_addra_77[8:0];
  assign weightRam_4_13_dina = sData_payload;
  assign weightRam_4_14_wea = weav_4_14;
  assign weightRam_4_14_addrb = weightRead_4_addr;
  assign weightData_4_14 = weightRam_4_14_doutb;
  assign weightRam_4_14_addra = _zz_addra_78[8:0];
  assign weightRam_4_14_dina = sData_payload;
  assign weightRam_4_15_wea = weav_4_15;
  assign weightRam_4_15_addrb = weightRead_4_addr;
  assign weightData_4_15 = weightRam_4_15_doutb;
  assign weightRam_4_15_addra = _zz_addra_79[8:0];
  assign weightRam_4_15_dina = sData_payload;
  assign weightRam_5_0_wea = weav_5_0;
  assign weightRam_5_0_addrb = weightRead_5_addr;
  assign weightData_5_0 = weightRam_5_0_doutb;
  assign weightRam_5_0_addra = _zz_addra_80[8:0];
  assign weightRam_5_0_dina = sData_payload;
  assign weightRam_5_1_wea = weav_5_1;
  assign weightRam_5_1_addrb = weightRead_5_addr;
  assign weightData_5_1 = weightRam_5_1_doutb;
  assign weightRam_5_1_addra = _zz_addra_81[8:0];
  assign weightRam_5_1_dina = sData_payload;
  assign weightRam_5_2_wea = weav_5_2;
  assign weightRam_5_2_addrb = weightRead_5_addr;
  assign weightData_5_2 = weightRam_5_2_doutb;
  assign weightRam_5_2_addra = _zz_addra_82[8:0];
  assign weightRam_5_2_dina = sData_payload;
  assign weightRam_5_3_wea = weav_5_3;
  assign weightRam_5_3_addrb = weightRead_5_addr;
  assign weightData_5_3 = weightRam_5_3_doutb;
  assign weightRam_5_3_addra = _zz_addra_83[8:0];
  assign weightRam_5_3_dina = sData_payload;
  assign weightRam_5_4_wea = weav_5_4;
  assign weightRam_5_4_addrb = weightRead_5_addr;
  assign weightData_5_4 = weightRam_5_4_doutb;
  assign weightRam_5_4_addra = _zz_addra_84[8:0];
  assign weightRam_5_4_dina = sData_payload;
  assign weightRam_5_5_wea = weav_5_5;
  assign weightRam_5_5_addrb = weightRead_5_addr;
  assign weightData_5_5 = weightRam_5_5_doutb;
  assign weightRam_5_5_addra = _zz_addra_85[8:0];
  assign weightRam_5_5_dina = sData_payload;
  assign weightRam_5_6_wea = weav_5_6;
  assign weightRam_5_6_addrb = weightRead_5_addr;
  assign weightData_5_6 = weightRam_5_6_doutb;
  assign weightRam_5_6_addra = _zz_addra_86[8:0];
  assign weightRam_5_6_dina = sData_payload;
  assign weightRam_5_7_wea = weav_5_7;
  assign weightRam_5_7_addrb = weightRead_5_addr;
  assign weightData_5_7 = weightRam_5_7_doutb;
  assign weightRam_5_7_addra = _zz_addra_87[8:0];
  assign weightRam_5_7_dina = sData_payload;
  assign weightRam_5_8_wea = weav_5_8;
  assign weightRam_5_8_addrb = weightRead_5_addr;
  assign weightData_5_8 = weightRam_5_8_doutb;
  assign weightRam_5_8_addra = _zz_addra_88[8:0];
  assign weightRam_5_8_dina = sData_payload;
  assign weightRam_5_9_wea = weav_5_9;
  assign weightRam_5_9_addrb = weightRead_5_addr;
  assign weightData_5_9 = weightRam_5_9_doutb;
  assign weightRam_5_9_addra = _zz_addra_89[8:0];
  assign weightRam_5_9_dina = sData_payload;
  assign weightRam_5_10_wea = weav_5_10;
  assign weightRam_5_10_addrb = weightRead_5_addr;
  assign weightData_5_10 = weightRam_5_10_doutb;
  assign weightRam_5_10_addra = _zz_addra_90[8:0];
  assign weightRam_5_10_dina = sData_payload;
  assign weightRam_5_11_wea = weav_5_11;
  assign weightRam_5_11_addrb = weightRead_5_addr;
  assign weightData_5_11 = weightRam_5_11_doutb;
  assign weightRam_5_11_addra = _zz_addra_91[8:0];
  assign weightRam_5_11_dina = sData_payload;
  assign weightRam_5_12_wea = weav_5_12;
  assign weightRam_5_12_addrb = weightRead_5_addr;
  assign weightData_5_12 = weightRam_5_12_doutb;
  assign weightRam_5_12_addra = _zz_addra_92[8:0];
  assign weightRam_5_12_dina = sData_payload;
  assign weightRam_5_13_wea = weav_5_13;
  assign weightRam_5_13_addrb = weightRead_5_addr;
  assign weightData_5_13 = weightRam_5_13_doutb;
  assign weightRam_5_13_addra = _zz_addra_93[8:0];
  assign weightRam_5_13_dina = sData_payload;
  assign weightRam_5_14_wea = weav_5_14;
  assign weightRam_5_14_addrb = weightRead_5_addr;
  assign weightData_5_14 = weightRam_5_14_doutb;
  assign weightRam_5_14_addra = _zz_addra_94[8:0];
  assign weightRam_5_14_dina = sData_payload;
  assign weightRam_5_15_wea = weav_5_15;
  assign weightRam_5_15_addrb = weightRead_5_addr;
  assign weightData_5_15 = weightRam_5_15_doutb;
  assign weightRam_5_15_addra = _zz_addra_95[8:0];
  assign weightRam_5_15_dina = sData_payload;
  assign weightRam_6_0_wea = weav_6_0;
  assign weightRam_6_0_addrb = weightRead_6_addr;
  assign weightData_6_0 = weightRam_6_0_doutb;
  assign weightRam_6_0_addra = _zz_addra_96[8:0];
  assign weightRam_6_0_dina = sData_payload;
  assign weightRam_6_1_wea = weav_6_1;
  assign weightRam_6_1_addrb = weightRead_6_addr;
  assign weightData_6_1 = weightRam_6_1_doutb;
  assign weightRam_6_1_addra = _zz_addra_97[8:0];
  assign weightRam_6_1_dina = sData_payload;
  assign weightRam_6_2_wea = weav_6_2;
  assign weightRam_6_2_addrb = weightRead_6_addr;
  assign weightData_6_2 = weightRam_6_2_doutb;
  assign weightRam_6_2_addra = _zz_addra_98[8:0];
  assign weightRam_6_2_dina = sData_payload;
  assign weightRam_6_3_wea = weav_6_3;
  assign weightRam_6_3_addrb = weightRead_6_addr;
  assign weightData_6_3 = weightRam_6_3_doutb;
  assign weightRam_6_3_addra = _zz_addra_99[8:0];
  assign weightRam_6_3_dina = sData_payload;
  assign weightRam_6_4_wea = weav_6_4;
  assign weightRam_6_4_addrb = weightRead_6_addr;
  assign weightData_6_4 = weightRam_6_4_doutb;
  assign weightRam_6_4_addra = _zz_addra_100[8:0];
  assign weightRam_6_4_dina = sData_payload;
  assign weightRam_6_5_wea = weav_6_5;
  assign weightRam_6_5_addrb = weightRead_6_addr;
  assign weightData_6_5 = weightRam_6_5_doutb;
  assign weightRam_6_5_addra = _zz_addra_101[8:0];
  assign weightRam_6_5_dina = sData_payload;
  assign weightRam_6_6_wea = weav_6_6;
  assign weightRam_6_6_addrb = weightRead_6_addr;
  assign weightData_6_6 = weightRam_6_6_doutb;
  assign weightRam_6_6_addra = _zz_addra_102[8:0];
  assign weightRam_6_6_dina = sData_payload;
  assign weightRam_6_7_wea = weav_6_7;
  assign weightRam_6_7_addrb = weightRead_6_addr;
  assign weightData_6_7 = weightRam_6_7_doutb;
  assign weightRam_6_7_addra = _zz_addra_103[8:0];
  assign weightRam_6_7_dina = sData_payload;
  assign weightRam_6_8_wea = weav_6_8;
  assign weightRam_6_8_addrb = weightRead_6_addr;
  assign weightData_6_8 = weightRam_6_8_doutb;
  assign weightRam_6_8_addra = _zz_addra_104[8:0];
  assign weightRam_6_8_dina = sData_payload;
  assign weightRam_6_9_wea = weav_6_9;
  assign weightRam_6_9_addrb = weightRead_6_addr;
  assign weightData_6_9 = weightRam_6_9_doutb;
  assign weightRam_6_9_addra = _zz_addra_105[8:0];
  assign weightRam_6_9_dina = sData_payload;
  assign weightRam_6_10_wea = weav_6_10;
  assign weightRam_6_10_addrb = weightRead_6_addr;
  assign weightData_6_10 = weightRam_6_10_doutb;
  assign weightRam_6_10_addra = _zz_addra_106[8:0];
  assign weightRam_6_10_dina = sData_payload;
  assign weightRam_6_11_wea = weav_6_11;
  assign weightRam_6_11_addrb = weightRead_6_addr;
  assign weightData_6_11 = weightRam_6_11_doutb;
  assign weightRam_6_11_addra = _zz_addra_107[8:0];
  assign weightRam_6_11_dina = sData_payload;
  assign weightRam_6_12_wea = weav_6_12;
  assign weightRam_6_12_addrb = weightRead_6_addr;
  assign weightData_6_12 = weightRam_6_12_doutb;
  assign weightRam_6_12_addra = _zz_addra_108[8:0];
  assign weightRam_6_12_dina = sData_payload;
  assign weightRam_6_13_wea = weav_6_13;
  assign weightRam_6_13_addrb = weightRead_6_addr;
  assign weightData_6_13 = weightRam_6_13_doutb;
  assign weightRam_6_13_addra = _zz_addra_109[8:0];
  assign weightRam_6_13_dina = sData_payload;
  assign weightRam_6_14_wea = weav_6_14;
  assign weightRam_6_14_addrb = weightRead_6_addr;
  assign weightData_6_14 = weightRam_6_14_doutb;
  assign weightRam_6_14_addra = _zz_addra_110[8:0];
  assign weightRam_6_14_dina = sData_payload;
  assign weightRam_6_15_wea = weav_6_15;
  assign weightRam_6_15_addrb = weightRead_6_addr;
  assign weightData_6_15 = weightRam_6_15_doutb;
  assign weightRam_6_15_addra = _zz_addra_111[8:0];
  assign weightRam_6_15_dina = sData_payload;
  assign weightRam_7_0_wea = weav_7_0;
  assign weightRam_7_0_addrb = weightRead_7_addr;
  assign weightData_7_0 = weightRam_7_0_doutb;
  assign weightRam_7_0_addra = _zz_addra_112[8:0];
  assign weightRam_7_0_dina = sData_payload;
  assign weightRam_7_1_wea = weav_7_1;
  assign weightRam_7_1_addrb = weightRead_7_addr;
  assign weightData_7_1 = weightRam_7_1_doutb;
  assign weightRam_7_1_addra = _zz_addra_113[8:0];
  assign weightRam_7_1_dina = sData_payload;
  assign weightRam_7_2_wea = weav_7_2;
  assign weightRam_7_2_addrb = weightRead_7_addr;
  assign weightData_7_2 = weightRam_7_2_doutb;
  assign weightRam_7_2_addra = _zz_addra_114[8:0];
  assign weightRam_7_2_dina = sData_payload;
  assign weightRam_7_3_wea = weav_7_3;
  assign weightRam_7_3_addrb = weightRead_7_addr;
  assign weightData_7_3 = weightRam_7_3_doutb;
  assign weightRam_7_3_addra = _zz_addra_115[8:0];
  assign weightRam_7_3_dina = sData_payload;
  assign weightRam_7_4_wea = weav_7_4;
  assign weightRam_7_4_addrb = weightRead_7_addr;
  assign weightData_7_4 = weightRam_7_4_doutb;
  assign weightRam_7_4_addra = _zz_addra_116[8:0];
  assign weightRam_7_4_dina = sData_payload;
  assign weightRam_7_5_wea = weav_7_5;
  assign weightRam_7_5_addrb = weightRead_7_addr;
  assign weightData_7_5 = weightRam_7_5_doutb;
  assign weightRam_7_5_addra = _zz_addra_117[8:0];
  assign weightRam_7_5_dina = sData_payload;
  assign weightRam_7_6_wea = weav_7_6;
  assign weightRam_7_6_addrb = weightRead_7_addr;
  assign weightData_7_6 = weightRam_7_6_doutb;
  assign weightRam_7_6_addra = _zz_addra_118[8:0];
  assign weightRam_7_6_dina = sData_payload;
  assign weightRam_7_7_wea = weav_7_7;
  assign weightRam_7_7_addrb = weightRead_7_addr;
  assign weightData_7_7 = weightRam_7_7_doutb;
  assign weightRam_7_7_addra = _zz_addra_119[8:0];
  assign weightRam_7_7_dina = sData_payload;
  assign weightRam_7_8_wea = weav_7_8;
  assign weightRam_7_8_addrb = weightRead_7_addr;
  assign weightData_7_8 = weightRam_7_8_doutb;
  assign weightRam_7_8_addra = _zz_addra_120[8:0];
  assign weightRam_7_8_dina = sData_payload;
  assign weightRam_7_9_wea = weav_7_9;
  assign weightRam_7_9_addrb = weightRead_7_addr;
  assign weightData_7_9 = weightRam_7_9_doutb;
  assign weightRam_7_9_addra = _zz_addra_121[8:0];
  assign weightRam_7_9_dina = sData_payload;
  assign weightRam_7_10_wea = weav_7_10;
  assign weightRam_7_10_addrb = weightRead_7_addr;
  assign weightData_7_10 = weightRam_7_10_doutb;
  assign weightRam_7_10_addra = _zz_addra_122[8:0];
  assign weightRam_7_10_dina = sData_payload;
  assign weightRam_7_11_wea = weav_7_11;
  assign weightRam_7_11_addrb = weightRead_7_addr;
  assign weightData_7_11 = weightRam_7_11_doutb;
  assign weightRam_7_11_addra = _zz_addra_123[8:0];
  assign weightRam_7_11_dina = sData_payload;
  assign weightRam_7_12_wea = weav_7_12;
  assign weightRam_7_12_addrb = weightRead_7_addr;
  assign weightData_7_12 = weightRam_7_12_doutb;
  assign weightRam_7_12_addra = _zz_addra_124[8:0];
  assign weightRam_7_12_dina = sData_payload;
  assign weightRam_7_13_wea = weav_7_13;
  assign weightRam_7_13_addrb = weightRead_7_addr;
  assign weightData_7_13 = weightRam_7_13_doutb;
  assign weightRam_7_13_addra = _zz_addra_125[8:0];
  assign weightRam_7_13_dina = sData_payload;
  assign weightRam_7_14_wea = weav_7_14;
  assign weightRam_7_14_addrb = weightRead_7_addr;
  assign weightData_7_14 = weightRam_7_14_doutb;
  assign weightRam_7_14_addra = _zz_addra_126[8:0];
  assign weightRam_7_14_dina = sData_payload;
  assign weightRam_7_15_wea = weav_7_15;
  assign weightRam_7_15_addrb = weightRead_7_addr;
  assign weightData_7_15 = weightRam_7_15_doutb;
  assign weightRam_7_15_addra = _zz_addra_127[8:0];
  assign weightRam_7_15_dina = sData_payload;
  assign weightRam_8_0_wea = weav_8_0;
  assign weightRam_8_0_addrb = weightRead_8_addr;
  assign weightData_8_0 = weightRam_8_0_doutb;
  assign weightRam_8_0_addra = _zz_addra_128[8:0];
  assign weightRam_8_0_dina = sData_payload;
  assign weightRam_8_1_wea = weav_8_1;
  assign weightRam_8_1_addrb = weightRead_8_addr;
  assign weightData_8_1 = weightRam_8_1_doutb;
  assign weightRam_8_1_addra = _zz_addra_129[8:0];
  assign weightRam_8_1_dina = sData_payload;
  assign weightRam_8_2_wea = weav_8_2;
  assign weightRam_8_2_addrb = weightRead_8_addr;
  assign weightData_8_2 = weightRam_8_2_doutb;
  assign weightRam_8_2_addra = _zz_addra_130[8:0];
  assign weightRam_8_2_dina = sData_payload;
  assign weightRam_8_3_wea = weav_8_3;
  assign weightRam_8_3_addrb = weightRead_8_addr;
  assign weightData_8_3 = weightRam_8_3_doutb;
  assign weightRam_8_3_addra = _zz_addra_131[8:0];
  assign weightRam_8_3_dina = sData_payload;
  assign weightRam_8_4_wea = weav_8_4;
  assign weightRam_8_4_addrb = weightRead_8_addr;
  assign weightData_8_4 = weightRam_8_4_doutb;
  assign weightRam_8_4_addra = _zz_addra_132[8:0];
  assign weightRam_8_4_dina = sData_payload;
  assign weightRam_8_5_wea = weav_8_5;
  assign weightRam_8_5_addrb = weightRead_8_addr;
  assign weightData_8_5 = weightRam_8_5_doutb;
  assign weightRam_8_5_addra = _zz_addra_133[8:0];
  assign weightRam_8_5_dina = sData_payload;
  assign weightRam_8_6_wea = weav_8_6;
  assign weightRam_8_6_addrb = weightRead_8_addr;
  assign weightData_8_6 = weightRam_8_6_doutb;
  assign weightRam_8_6_addra = _zz_addra_134[8:0];
  assign weightRam_8_6_dina = sData_payload;
  assign weightRam_8_7_wea = weav_8_7;
  assign weightRam_8_7_addrb = weightRead_8_addr;
  assign weightData_8_7 = weightRam_8_7_doutb;
  assign weightRam_8_7_addra = _zz_addra_135[8:0];
  assign weightRam_8_7_dina = sData_payload;
  assign weightRam_8_8_wea = weav_8_8;
  assign weightRam_8_8_addrb = weightRead_8_addr;
  assign weightData_8_8 = weightRam_8_8_doutb;
  assign weightRam_8_8_addra = _zz_addra_136[8:0];
  assign weightRam_8_8_dina = sData_payload;
  assign weightRam_8_9_wea = weav_8_9;
  assign weightRam_8_9_addrb = weightRead_8_addr;
  assign weightData_8_9 = weightRam_8_9_doutb;
  assign weightRam_8_9_addra = _zz_addra_137[8:0];
  assign weightRam_8_9_dina = sData_payload;
  assign weightRam_8_10_wea = weav_8_10;
  assign weightRam_8_10_addrb = weightRead_8_addr;
  assign weightData_8_10 = weightRam_8_10_doutb;
  assign weightRam_8_10_addra = _zz_addra_138[8:0];
  assign weightRam_8_10_dina = sData_payload;
  assign weightRam_8_11_wea = weav_8_11;
  assign weightRam_8_11_addrb = weightRead_8_addr;
  assign weightData_8_11 = weightRam_8_11_doutb;
  assign weightRam_8_11_addra = _zz_addra_139[8:0];
  assign weightRam_8_11_dina = sData_payload;
  assign weightRam_8_12_wea = weav_8_12;
  assign weightRam_8_12_addrb = weightRead_8_addr;
  assign weightData_8_12 = weightRam_8_12_doutb;
  assign weightRam_8_12_addra = _zz_addra_140[8:0];
  assign weightRam_8_12_dina = sData_payload;
  assign weightRam_8_13_wea = weav_8_13;
  assign weightRam_8_13_addrb = weightRead_8_addr;
  assign weightData_8_13 = weightRam_8_13_doutb;
  assign weightRam_8_13_addra = _zz_addra_141[8:0];
  assign weightRam_8_13_dina = sData_payload;
  assign weightRam_8_14_wea = weav_8_14;
  assign weightRam_8_14_addrb = weightRead_8_addr;
  assign weightData_8_14 = weightRam_8_14_doutb;
  assign weightRam_8_14_addra = _zz_addra_142[8:0];
  assign weightRam_8_14_dina = sData_payload;
  assign weightRam_8_15_wea = weav_8_15;
  assign weightRam_8_15_addrb = weightRead_8_addr;
  assign weightData_8_15 = weightRam_8_15_doutb;
  assign weightRam_8_15_addra = _zz_addra_143[8:0];
  assign weightRam_8_15_dina = sData_payload;
  assign sData_fire_4 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_4 = (((fsm_currentState & LoadWeightEnum_COPY_BIAS) != 6'b000000) && sData_fire_4);
  assign sData_fire_5 = (sData_valid && sData_ready);
  assign when_WaCounter_l12_7 = (copyBias_copyCnt_count == _zz_when_WaCounter_l12_7);
  always @(*) begin
    if(when_WaCounter_l12_7) begin
      copyBias_copyCnt_valid = 1'b1;
    end else begin
      copyBias_copyCnt_valid = 1'b0;
    end
  end

  assign copyBias_ram_wea = (((fsm_currentState & LoadWeightEnum_COPY_BIAS) != 6'b000000) && sData_fire_5);
  assign copyBias_ram_dina = sData_payload;
  assign copyBias_ram_addra = copyBias_copyCnt_count;
  assign copyBias_ram_addrb = biasRead_addr;
  assign biasRead_data = copyBias_ram_doutb;
  assign fsm_copyBiasEnd = copyBias_copyCnt_valid;
  assign sData_fire_6 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_5 = (((fsm_currentState & LoadWeightEnum_COPY_SCALE) != 6'b000000) && sData_fire_6);
  assign sData_fire_7 = (sData_valid && sData_ready);
  assign when_WaCounter_l12_8 = (copyScale_copyCnt_count == _zz_when_WaCounter_l12_8);
  always @(*) begin
    if(when_WaCounter_l12_8) begin
      copyScale_copyCnt_valid = 1'b1;
    end else begin
      copyScale_copyCnt_valid = 1'b0;
    end
  end

  assign copyScale_ram_wea = (((fsm_currentState & LoadWeightEnum_COPY_SCALE) != 6'b000000) && sData_fire_7);
  assign copyScale_ram_dina = sData_payload;
  assign copyScale_ram_addra = copyScale_copyCnt_count;
  assign copyScale_ram_addrb = scaleRead_addr;
  assign scaleRead_data = copyScale_ram_doutb;
  assign fsm_copyScaleEnd = copyScale_copyCnt_valid;
  assign sData_fire_8 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_6 = (((fsm_currentState & LoadWeightEnum_COPY_SHIFT) != 6'b000000) && sData_fire_8);
  assign sData_fire_9 = (sData_valid && sData_ready);
  assign when_WaCounter_l12_9 = (copyShift_copyCnt_count == _zz_when_WaCounter_l12_9);
  always @(*) begin
    if(when_WaCounter_l12_9) begin
      copyShift_copyCnt_valid = 1'b1;
    end else begin
      copyShift_copyCnt_valid = 1'b0;
    end
  end

  assign copyShift_ram_wea = (((fsm_currentState & LoadWeightEnum_COPY_SHIFT) != 6'b000000) && sData_fire_9);
  assign copyShift_ram_dina = sData_payload;
  assign copyShift_ram_addra = copyShift_copyCnt_count;
  assign copyShift_ram_addrb = shiftRead_addr;
  assign shiftRead_data = copyShift_ram_doutb;
  assign fsm_copyShiftEnd = copyShift_copyCnt_valid;
  assign when_WaUtil_l29 = (((fsm_currentState & LoadWeightEnum_COPY_SHIFT) != 6'b000000) && ((fsm_nextState & LoadWeightEnum_IDLE) != 6'b000000));
  always @(*) begin
    if(when_WaUtil_l29) begin
      copyWeightDone = 1'b1;
    end else begin
      copyWeightDone = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      fsm_currentState <= LoadWeightEnum_IDLE;
      init_count <= 3'b000;
      copyWeightCnt_count <= 13'h0;
      copyWeightTimes_count <= 4'b0000;
      channelInCnt_count <= 8'h0;
      computeChannelOut_count <= 4'b0000;
      times_count <= 4'b0000;
      channelOutCnt_count <= 12'h0;
      addr_0_0 <= 13'h0;
      addr_0_1 <= 13'h0;
      addr_0_2 <= 13'h0;
      addr_0_3 <= 13'h0;
      addr_0_4 <= 13'h0;
      addr_0_5 <= 13'h0;
      addr_0_6 <= 13'h0;
      addr_0_7 <= 13'h0;
      addr_0_8 <= 13'h0;
      addr_0_9 <= 13'h0;
      addr_0_10 <= 13'h0;
      addr_0_11 <= 13'h0;
      addr_0_12 <= 13'h0;
      addr_0_13 <= 13'h0;
      addr_0_14 <= 13'h0;
      addr_0_15 <= 13'h0;
      addr_1_0 <= 13'h0;
      addr_1_1 <= 13'h0;
      addr_1_2 <= 13'h0;
      addr_1_3 <= 13'h0;
      addr_1_4 <= 13'h0;
      addr_1_5 <= 13'h0;
      addr_1_6 <= 13'h0;
      addr_1_7 <= 13'h0;
      addr_1_8 <= 13'h0;
      addr_1_9 <= 13'h0;
      addr_1_10 <= 13'h0;
      addr_1_11 <= 13'h0;
      addr_1_12 <= 13'h0;
      addr_1_13 <= 13'h0;
      addr_1_14 <= 13'h0;
      addr_1_15 <= 13'h0;
      addr_2_0 <= 13'h0;
      addr_2_1 <= 13'h0;
      addr_2_2 <= 13'h0;
      addr_2_3 <= 13'h0;
      addr_2_4 <= 13'h0;
      addr_2_5 <= 13'h0;
      addr_2_6 <= 13'h0;
      addr_2_7 <= 13'h0;
      addr_2_8 <= 13'h0;
      addr_2_9 <= 13'h0;
      addr_2_10 <= 13'h0;
      addr_2_11 <= 13'h0;
      addr_2_12 <= 13'h0;
      addr_2_13 <= 13'h0;
      addr_2_14 <= 13'h0;
      addr_2_15 <= 13'h0;
      addr_3_0 <= 13'h0;
      addr_3_1 <= 13'h0;
      addr_3_2 <= 13'h0;
      addr_3_3 <= 13'h0;
      addr_3_4 <= 13'h0;
      addr_3_5 <= 13'h0;
      addr_3_6 <= 13'h0;
      addr_3_7 <= 13'h0;
      addr_3_8 <= 13'h0;
      addr_3_9 <= 13'h0;
      addr_3_10 <= 13'h0;
      addr_3_11 <= 13'h0;
      addr_3_12 <= 13'h0;
      addr_3_13 <= 13'h0;
      addr_3_14 <= 13'h0;
      addr_3_15 <= 13'h0;
      addr_4_0 <= 13'h0;
      addr_4_1 <= 13'h0;
      addr_4_2 <= 13'h0;
      addr_4_3 <= 13'h0;
      addr_4_4 <= 13'h0;
      addr_4_5 <= 13'h0;
      addr_4_6 <= 13'h0;
      addr_4_7 <= 13'h0;
      addr_4_8 <= 13'h0;
      addr_4_9 <= 13'h0;
      addr_4_10 <= 13'h0;
      addr_4_11 <= 13'h0;
      addr_4_12 <= 13'h0;
      addr_4_13 <= 13'h0;
      addr_4_14 <= 13'h0;
      addr_4_15 <= 13'h0;
      addr_5_0 <= 13'h0;
      addr_5_1 <= 13'h0;
      addr_5_2 <= 13'h0;
      addr_5_3 <= 13'h0;
      addr_5_4 <= 13'h0;
      addr_5_5 <= 13'h0;
      addr_5_6 <= 13'h0;
      addr_5_7 <= 13'h0;
      addr_5_8 <= 13'h0;
      addr_5_9 <= 13'h0;
      addr_5_10 <= 13'h0;
      addr_5_11 <= 13'h0;
      addr_5_12 <= 13'h0;
      addr_5_13 <= 13'h0;
      addr_5_14 <= 13'h0;
      addr_5_15 <= 13'h0;
      addr_6_0 <= 13'h0;
      addr_6_1 <= 13'h0;
      addr_6_2 <= 13'h0;
      addr_6_3 <= 13'h0;
      addr_6_4 <= 13'h0;
      addr_6_5 <= 13'h0;
      addr_6_6 <= 13'h0;
      addr_6_7 <= 13'h0;
      addr_6_8 <= 13'h0;
      addr_6_9 <= 13'h0;
      addr_6_10 <= 13'h0;
      addr_6_11 <= 13'h0;
      addr_6_12 <= 13'h0;
      addr_6_13 <= 13'h0;
      addr_6_14 <= 13'h0;
      addr_6_15 <= 13'h0;
      addr_7_0 <= 13'h0;
      addr_7_1 <= 13'h0;
      addr_7_2 <= 13'h0;
      addr_7_3 <= 13'h0;
      addr_7_4 <= 13'h0;
      addr_7_5 <= 13'h0;
      addr_7_6 <= 13'h0;
      addr_7_7 <= 13'h0;
      addr_7_8 <= 13'h0;
      addr_7_9 <= 13'h0;
      addr_7_10 <= 13'h0;
      addr_7_11 <= 13'h0;
      addr_7_12 <= 13'h0;
      addr_7_13 <= 13'h0;
      addr_7_14 <= 13'h0;
      addr_7_15 <= 13'h0;
      addr_8_0 <= 13'h0;
      addr_8_1 <= 13'h0;
      addr_8_2 <= 13'h0;
      addr_8_3 <= 13'h0;
      addr_8_4 <= 13'h0;
      addr_8_5 <= 13'h0;
      addr_8_6 <= 13'h0;
      addr_8_7 <= 13'h0;
      addr_8_8 <= 13'h0;
      addr_8_9 <= 13'h0;
      addr_8_10 <= 13'h0;
      addr_8_11 <= 13'h0;
      addr_8_12 <= 13'h0;
      addr_8_13 <= 13'h0;
      addr_8_14 <= 13'h0;
      addr_8_15 <= 13'h0;
      copyBias_copyCnt_count <= 8'h0;
      copyScale_copyCnt_count <= 8'h0;
      copyShift_copyCnt_count <= 8'h0;
    end else begin
      if(softReset) begin
      fsm_currentState <= LoadWeightEnum_IDLE;
      init_count <= 3'b000;
      copyWeightCnt_count <= 13'h0;
      copyWeightTimes_count <= 4'b0000;
      channelInCnt_count <= 8'h0;
      computeChannelOut_count <= 4'b0000;
      times_count <= 4'b0000;
      channelOutCnt_count <= 12'h0;
      addr_0_0 <= 13'h0;
      addr_0_1 <= 13'h0;
      addr_0_2 <= 13'h0;
      addr_0_3 <= 13'h0;
      addr_0_4 <= 13'h0;
      addr_0_5 <= 13'h0;
      addr_0_6 <= 13'h0;
      addr_0_7 <= 13'h0;
      addr_0_8 <= 13'h0;
      addr_0_9 <= 13'h0;
      addr_0_10 <= 13'h0;
      addr_0_11 <= 13'h0;
      addr_0_12 <= 13'h0;
      addr_0_13 <= 13'h0;
      addr_0_14 <= 13'h0;
      addr_0_15 <= 13'h0;
      addr_1_0 <= 13'h0;
      addr_1_1 <= 13'h0;
      addr_1_2 <= 13'h0;
      addr_1_3 <= 13'h0;
      addr_1_4 <= 13'h0;
      addr_1_5 <= 13'h0;
      addr_1_6 <= 13'h0;
      addr_1_7 <= 13'h0;
      addr_1_8 <= 13'h0;
      addr_1_9 <= 13'h0;
      addr_1_10 <= 13'h0;
      addr_1_11 <= 13'h0;
      addr_1_12 <= 13'h0;
      addr_1_13 <= 13'h0;
      addr_1_14 <= 13'h0;
      addr_1_15 <= 13'h0;
      addr_2_0 <= 13'h0;
      addr_2_1 <= 13'h0;
      addr_2_2 <= 13'h0;
      addr_2_3 <= 13'h0;
      addr_2_4 <= 13'h0;
      addr_2_5 <= 13'h0;
      addr_2_6 <= 13'h0;
      addr_2_7 <= 13'h0;
      addr_2_8 <= 13'h0;
      addr_2_9 <= 13'h0;
      addr_2_10 <= 13'h0;
      addr_2_11 <= 13'h0;
      addr_2_12 <= 13'h0;
      addr_2_13 <= 13'h0;
      addr_2_14 <= 13'h0;
      addr_2_15 <= 13'h0;
      addr_3_0 <= 13'h0;
      addr_3_1 <= 13'h0;
      addr_3_2 <= 13'h0;
      addr_3_3 <= 13'h0;
      addr_3_4 <= 13'h0;
      addr_3_5 <= 13'h0;
      addr_3_6 <= 13'h0;
      addr_3_7 <= 13'h0;
      addr_3_8 <= 13'h0;
      addr_3_9 <= 13'h0;
      addr_3_10 <= 13'h0;
      addr_3_11 <= 13'h0;
      addr_3_12 <= 13'h0;
      addr_3_13 <= 13'h0;
      addr_3_14 <= 13'h0;
      addr_3_15 <= 13'h0;
      addr_4_0 <= 13'h0;
      addr_4_1 <= 13'h0;
      addr_4_2 <= 13'h0;
      addr_4_3 <= 13'h0;
      addr_4_4 <= 13'h0;
      addr_4_5 <= 13'h0;
      addr_4_6 <= 13'h0;
      addr_4_7 <= 13'h0;
      addr_4_8 <= 13'h0;
      addr_4_9 <= 13'h0;
      addr_4_10 <= 13'h0;
      addr_4_11 <= 13'h0;
      addr_4_12 <= 13'h0;
      addr_4_13 <= 13'h0;
      addr_4_14 <= 13'h0;
      addr_4_15 <= 13'h0;
      addr_5_0 <= 13'h0;
      addr_5_1 <= 13'h0;
      addr_5_2 <= 13'h0;
      addr_5_3 <= 13'h0;
      addr_5_4 <= 13'h0;
      addr_5_5 <= 13'h0;
      addr_5_6 <= 13'h0;
      addr_5_7 <= 13'h0;
      addr_5_8 <= 13'h0;
      addr_5_9 <= 13'h0;
      addr_5_10 <= 13'h0;
      addr_5_11 <= 13'h0;
      addr_5_12 <= 13'h0;
      addr_5_13 <= 13'h0;
      addr_5_14 <= 13'h0;
      addr_5_15 <= 13'h0;
      addr_6_0 <= 13'h0;
      addr_6_1 <= 13'h0;
      addr_6_2 <= 13'h0;
      addr_6_3 <= 13'h0;
      addr_6_4 <= 13'h0;
      addr_6_5 <= 13'h0;
      addr_6_6 <= 13'h0;
      addr_6_7 <= 13'h0;
      addr_6_8 <= 13'h0;
      addr_6_9 <= 13'h0;
      addr_6_10 <= 13'h0;
      addr_6_11 <= 13'h0;
      addr_6_12 <= 13'h0;
      addr_6_13 <= 13'h0;
      addr_6_14 <= 13'h0;
      addr_6_15 <= 13'h0;
      addr_7_0 <= 13'h0;
      addr_7_1 <= 13'h0;
      addr_7_2 <= 13'h0;
      addr_7_3 <= 13'h0;
      addr_7_4 <= 13'h0;
      addr_7_5 <= 13'h0;
      addr_7_6 <= 13'h0;
      addr_7_7 <= 13'h0;
      addr_7_8 <= 13'h0;
      addr_7_9 <= 13'h0;
      addr_7_10 <= 13'h0;
      addr_7_11 <= 13'h0;
      addr_7_12 <= 13'h0;
      addr_7_13 <= 13'h0;
      addr_7_14 <= 13'h0;
      addr_7_15 <= 13'h0;
      addr_8_0 <= 13'h0;
      addr_8_1 <= 13'h0;
      addr_8_2 <= 13'h0;
      addr_8_3 <= 13'h0;
      addr_8_4 <= 13'h0;
      addr_8_5 <= 13'h0;
      addr_8_6 <= 13'h0;
      addr_8_7 <= 13'h0;
      addr_8_8 <= 13'h0;
      addr_8_9 <= 13'h0;
      addr_8_10 <= 13'h0;
      addr_8_11 <= 13'h0;
      addr_8_12 <= 13'h0;
      addr_8_13 <= 13'h0;
      addr_8_14 <= 13'h0;
      addr_8_15 <= 13'h0;
      copyBias_copyCnt_count <= 8'h0;
      copyScale_copyCnt_count <= 8'h0;
      copyShift_copyCnt_count <= 8'h0;
      end else begin
        fsm_currentState <= fsm_nextState;
        if(when_WaCounter_l17) begin
          init_count <= (init_count + 3'b001);
          if(init_valid) begin
            init_count <= 3'b000;
          end
        end
        if(when_WaCounter_l17_1) begin
          copyWeightCnt_count <= (copyWeightCnt_count + 13'h0001);
          if(copyWeightCnt_valid) begin
            copyWeightCnt_count <= 13'h0;
          end
        end
        if(copyWeightCnt_valid) begin
          copyWeightTimes_count <= (copyWeightTimes_count + 4'b0001);
          if(copyWeightTimes_valid) begin
            copyWeightTimes_count <= 4'b0000;
          end
        end
        if(when_WaCounter_l17_2) begin
          channelInCnt_count <= (channelInCnt_count + 8'h01);
          if(channelInCnt_valid) begin
            channelInCnt_count <= 8'h0;
          end
        end
        if(when_WaCounter_l17_3) begin
          computeChannelOut_count <= (computeChannelOut_count + 4'b0001);
          if(computeChannelOut_valid) begin
            computeChannelOut_count <= 4'b0000;
          end
        end
        if(computeChannelOut_valid) begin
          times_count <= (times_count + 4'b0001);
          if(times_valid) begin
            times_count <= 4'b0000;
          end
        end
        if(channelInCnt_valid) begin
          channelOutCnt_count <= (channelOutCnt_count + 12'h001);
          if(channelOutCnt_valid) begin
            channelOutCnt_count <= 12'h0;
          end
        end
        if(when_Weight_l250) begin
          channelInCnt_count <= 8'h0;
          computeChannelOut_count <= 4'b0000;
          times_count <= 4'b0000;
          channelOutCnt_count <= 12'h0;
        end
        if(weav_0_0) begin
          if(when_Weight_l326) begin
            addr_0_0 <= 13'h0;
          end else begin
            addr_0_0 <= (addr_0_0 + 13'h0001);
          end
        end
        if(weav_0_1) begin
          if(when_Weight_l326_1) begin
            addr_0_1 <= 13'h0;
          end else begin
            addr_0_1 <= (addr_0_1 + 13'h0001);
          end
        end
        if(weav_0_2) begin
          if(when_Weight_l326_2) begin
            addr_0_2 <= 13'h0;
          end else begin
            addr_0_2 <= (addr_0_2 + 13'h0001);
          end
        end
        if(weav_0_3) begin
          if(when_Weight_l326_3) begin
            addr_0_3 <= 13'h0;
          end else begin
            addr_0_3 <= (addr_0_3 + 13'h0001);
          end
        end
        if(weav_0_4) begin
          if(when_Weight_l326_4) begin
            addr_0_4 <= 13'h0;
          end else begin
            addr_0_4 <= (addr_0_4 + 13'h0001);
          end
        end
        if(weav_0_5) begin
          if(when_Weight_l326_5) begin
            addr_0_5 <= 13'h0;
          end else begin
            addr_0_5 <= (addr_0_5 + 13'h0001);
          end
        end
        if(weav_0_6) begin
          if(when_Weight_l326_6) begin
            addr_0_6 <= 13'h0;
          end else begin
            addr_0_6 <= (addr_0_6 + 13'h0001);
          end
        end
        if(weav_0_7) begin
          if(when_Weight_l326_7) begin
            addr_0_7 <= 13'h0;
          end else begin
            addr_0_7 <= (addr_0_7 + 13'h0001);
          end
        end
        if(weav_0_8) begin
          if(when_Weight_l326_8) begin
            addr_0_8 <= 13'h0;
          end else begin
            addr_0_8 <= (addr_0_8 + 13'h0001);
          end
        end
        if(weav_0_9) begin
          if(when_Weight_l326_9) begin
            addr_0_9 <= 13'h0;
          end else begin
            addr_0_9 <= (addr_0_9 + 13'h0001);
          end
        end
        if(weav_0_10) begin
          if(when_Weight_l326_10) begin
            addr_0_10 <= 13'h0;
          end else begin
            addr_0_10 <= (addr_0_10 + 13'h0001);
          end
        end
        if(weav_0_11) begin
          if(when_Weight_l326_11) begin
            addr_0_11 <= 13'h0;
          end else begin
            addr_0_11 <= (addr_0_11 + 13'h0001);
          end
        end
        if(weav_0_12) begin
          if(when_Weight_l326_12) begin
            addr_0_12 <= 13'h0;
          end else begin
            addr_0_12 <= (addr_0_12 + 13'h0001);
          end
        end
        if(weav_0_13) begin
          if(when_Weight_l326_13) begin
            addr_0_13 <= 13'h0;
          end else begin
            addr_0_13 <= (addr_0_13 + 13'h0001);
          end
        end
        if(weav_0_14) begin
          if(when_Weight_l326_14) begin
            addr_0_14 <= 13'h0;
          end else begin
            addr_0_14 <= (addr_0_14 + 13'h0001);
          end
        end
        if(weav_0_15) begin
          if(when_Weight_l326_15) begin
            addr_0_15 <= 13'h0;
          end else begin
            addr_0_15 <= (addr_0_15 + 13'h0001);
          end
        end
        if(weav_1_0) begin
          if(when_Weight_l326_16) begin
            addr_1_0 <= 13'h0;
          end else begin
            addr_1_0 <= (addr_1_0 + 13'h0001);
          end
        end
        if(weav_1_1) begin
          if(when_Weight_l326_17) begin
            addr_1_1 <= 13'h0;
          end else begin
            addr_1_1 <= (addr_1_1 + 13'h0001);
          end
        end
        if(weav_1_2) begin
          if(when_Weight_l326_18) begin
            addr_1_2 <= 13'h0;
          end else begin
            addr_1_2 <= (addr_1_2 + 13'h0001);
          end
        end
        if(weav_1_3) begin
          if(when_Weight_l326_19) begin
            addr_1_3 <= 13'h0;
          end else begin
            addr_1_3 <= (addr_1_3 + 13'h0001);
          end
        end
        if(weav_1_4) begin
          if(when_Weight_l326_20) begin
            addr_1_4 <= 13'h0;
          end else begin
            addr_1_4 <= (addr_1_4 + 13'h0001);
          end
        end
        if(weav_1_5) begin
          if(when_Weight_l326_21) begin
            addr_1_5 <= 13'h0;
          end else begin
            addr_1_5 <= (addr_1_5 + 13'h0001);
          end
        end
        if(weav_1_6) begin
          if(when_Weight_l326_22) begin
            addr_1_6 <= 13'h0;
          end else begin
            addr_1_6 <= (addr_1_6 + 13'h0001);
          end
        end
        if(weav_1_7) begin
          if(when_Weight_l326_23) begin
            addr_1_7 <= 13'h0;
          end else begin
            addr_1_7 <= (addr_1_7 + 13'h0001);
          end
        end
        if(weav_1_8) begin
          if(when_Weight_l326_24) begin
            addr_1_8 <= 13'h0;
          end else begin
            addr_1_8 <= (addr_1_8 + 13'h0001);
          end
        end
        if(weav_1_9) begin
          if(when_Weight_l326_25) begin
            addr_1_9 <= 13'h0;
          end else begin
            addr_1_9 <= (addr_1_9 + 13'h0001);
          end
        end
        if(weav_1_10) begin
          if(when_Weight_l326_26) begin
            addr_1_10 <= 13'h0;
          end else begin
            addr_1_10 <= (addr_1_10 + 13'h0001);
          end
        end
        if(weav_1_11) begin
          if(when_Weight_l326_27) begin
            addr_1_11 <= 13'h0;
          end else begin
            addr_1_11 <= (addr_1_11 + 13'h0001);
          end
        end
        if(weav_1_12) begin
          if(when_Weight_l326_28) begin
            addr_1_12 <= 13'h0;
          end else begin
            addr_1_12 <= (addr_1_12 + 13'h0001);
          end
        end
        if(weav_1_13) begin
          if(when_Weight_l326_29) begin
            addr_1_13 <= 13'h0;
          end else begin
            addr_1_13 <= (addr_1_13 + 13'h0001);
          end
        end
        if(weav_1_14) begin
          if(when_Weight_l326_30) begin
            addr_1_14 <= 13'h0;
          end else begin
            addr_1_14 <= (addr_1_14 + 13'h0001);
          end
        end
        if(weav_1_15) begin
          if(when_Weight_l326_31) begin
            addr_1_15 <= 13'h0;
          end else begin
            addr_1_15 <= (addr_1_15 + 13'h0001);
          end
        end
        if(weav_2_0) begin
          if(when_Weight_l326_32) begin
            addr_2_0 <= 13'h0;
          end else begin
            addr_2_0 <= (addr_2_0 + 13'h0001);
          end
        end
        if(weav_2_1) begin
          if(when_Weight_l326_33) begin
            addr_2_1 <= 13'h0;
          end else begin
            addr_2_1 <= (addr_2_1 + 13'h0001);
          end
        end
        if(weav_2_2) begin
          if(when_Weight_l326_34) begin
            addr_2_2 <= 13'h0;
          end else begin
            addr_2_2 <= (addr_2_2 + 13'h0001);
          end
        end
        if(weav_2_3) begin
          if(when_Weight_l326_35) begin
            addr_2_3 <= 13'h0;
          end else begin
            addr_2_3 <= (addr_2_3 + 13'h0001);
          end
        end
        if(weav_2_4) begin
          if(when_Weight_l326_36) begin
            addr_2_4 <= 13'h0;
          end else begin
            addr_2_4 <= (addr_2_4 + 13'h0001);
          end
        end
        if(weav_2_5) begin
          if(when_Weight_l326_37) begin
            addr_2_5 <= 13'h0;
          end else begin
            addr_2_5 <= (addr_2_5 + 13'h0001);
          end
        end
        if(weav_2_6) begin
          if(when_Weight_l326_38) begin
            addr_2_6 <= 13'h0;
          end else begin
            addr_2_6 <= (addr_2_6 + 13'h0001);
          end
        end
        if(weav_2_7) begin
          if(when_Weight_l326_39) begin
            addr_2_7 <= 13'h0;
          end else begin
            addr_2_7 <= (addr_2_7 + 13'h0001);
          end
        end
        if(weav_2_8) begin
          if(when_Weight_l326_40) begin
            addr_2_8 <= 13'h0;
          end else begin
            addr_2_8 <= (addr_2_8 + 13'h0001);
          end
        end
        if(weav_2_9) begin
          if(when_Weight_l326_41) begin
            addr_2_9 <= 13'h0;
          end else begin
            addr_2_9 <= (addr_2_9 + 13'h0001);
          end
        end
        if(weav_2_10) begin
          if(when_Weight_l326_42) begin
            addr_2_10 <= 13'h0;
          end else begin
            addr_2_10 <= (addr_2_10 + 13'h0001);
          end
        end
        if(weav_2_11) begin
          if(when_Weight_l326_43) begin
            addr_2_11 <= 13'h0;
          end else begin
            addr_2_11 <= (addr_2_11 + 13'h0001);
          end
        end
        if(weav_2_12) begin
          if(when_Weight_l326_44) begin
            addr_2_12 <= 13'h0;
          end else begin
            addr_2_12 <= (addr_2_12 + 13'h0001);
          end
        end
        if(weav_2_13) begin
          if(when_Weight_l326_45) begin
            addr_2_13 <= 13'h0;
          end else begin
            addr_2_13 <= (addr_2_13 + 13'h0001);
          end
        end
        if(weav_2_14) begin
          if(when_Weight_l326_46) begin
            addr_2_14 <= 13'h0;
          end else begin
            addr_2_14 <= (addr_2_14 + 13'h0001);
          end
        end
        if(weav_2_15) begin
          if(when_Weight_l326_47) begin
            addr_2_15 <= 13'h0;
          end else begin
            addr_2_15 <= (addr_2_15 + 13'h0001);
          end
        end
        if(weav_3_0) begin
          if(when_Weight_l326_48) begin
            addr_3_0 <= 13'h0;
          end else begin
            addr_3_0 <= (addr_3_0 + 13'h0001);
          end
        end
        if(weav_3_1) begin
          if(when_Weight_l326_49) begin
            addr_3_1 <= 13'h0;
          end else begin
            addr_3_1 <= (addr_3_1 + 13'h0001);
          end
        end
        if(weav_3_2) begin
          if(when_Weight_l326_50) begin
            addr_3_2 <= 13'h0;
          end else begin
            addr_3_2 <= (addr_3_2 + 13'h0001);
          end
        end
        if(weav_3_3) begin
          if(when_Weight_l326_51) begin
            addr_3_3 <= 13'h0;
          end else begin
            addr_3_3 <= (addr_3_3 + 13'h0001);
          end
        end
        if(weav_3_4) begin
          if(when_Weight_l326_52) begin
            addr_3_4 <= 13'h0;
          end else begin
            addr_3_4 <= (addr_3_4 + 13'h0001);
          end
        end
        if(weav_3_5) begin
          if(when_Weight_l326_53) begin
            addr_3_5 <= 13'h0;
          end else begin
            addr_3_5 <= (addr_3_5 + 13'h0001);
          end
        end
        if(weav_3_6) begin
          if(when_Weight_l326_54) begin
            addr_3_6 <= 13'h0;
          end else begin
            addr_3_6 <= (addr_3_6 + 13'h0001);
          end
        end
        if(weav_3_7) begin
          if(when_Weight_l326_55) begin
            addr_3_7 <= 13'h0;
          end else begin
            addr_3_7 <= (addr_3_7 + 13'h0001);
          end
        end
        if(weav_3_8) begin
          if(when_Weight_l326_56) begin
            addr_3_8 <= 13'h0;
          end else begin
            addr_3_8 <= (addr_3_8 + 13'h0001);
          end
        end
        if(weav_3_9) begin
          if(when_Weight_l326_57) begin
            addr_3_9 <= 13'h0;
          end else begin
            addr_3_9 <= (addr_3_9 + 13'h0001);
          end
        end
        if(weav_3_10) begin
          if(when_Weight_l326_58) begin
            addr_3_10 <= 13'h0;
          end else begin
            addr_3_10 <= (addr_3_10 + 13'h0001);
          end
        end
        if(weav_3_11) begin
          if(when_Weight_l326_59) begin
            addr_3_11 <= 13'h0;
          end else begin
            addr_3_11 <= (addr_3_11 + 13'h0001);
          end
        end
        if(weav_3_12) begin
          if(when_Weight_l326_60) begin
            addr_3_12 <= 13'h0;
          end else begin
            addr_3_12 <= (addr_3_12 + 13'h0001);
          end
        end
        if(weav_3_13) begin
          if(when_Weight_l326_61) begin
            addr_3_13 <= 13'h0;
          end else begin
            addr_3_13 <= (addr_3_13 + 13'h0001);
          end
        end
        if(weav_3_14) begin
          if(when_Weight_l326_62) begin
            addr_3_14 <= 13'h0;
          end else begin
            addr_3_14 <= (addr_3_14 + 13'h0001);
          end
        end
        if(weav_3_15) begin
          if(when_Weight_l326_63) begin
            addr_3_15 <= 13'h0;
          end else begin
            addr_3_15 <= (addr_3_15 + 13'h0001);
          end
        end
        if(weav_4_0) begin
          if(when_Weight_l326_64) begin
            addr_4_0 <= 13'h0;
          end else begin
            addr_4_0 <= (addr_4_0 + 13'h0001);
          end
        end
        if(weav_4_1) begin
          if(when_Weight_l326_65) begin
            addr_4_1 <= 13'h0;
          end else begin
            addr_4_1 <= (addr_4_1 + 13'h0001);
          end
        end
        if(weav_4_2) begin
          if(when_Weight_l326_66) begin
            addr_4_2 <= 13'h0;
          end else begin
            addr_4_2 <= (addr_4_2 + 13'h0001);
          end
        end
        if(weav_4_3) begin
          if(when_Weight_l326_67) begin
            addr_4_3 <= 13'h0;
          end else begin
            addr_4_3 <= (addr_4_3 + 13'h0001);
          end
        end
        if(weav_4_4) begin
          if(when_Weight_l326_68) begin
            addr_4_4 <= 13'h0;
          end else begin
            addr_4_4 <= (addr_4_4 + 13'h0001);
          end
        end
        if(weav_4_5) begin
          if(when_Weight_l326_69) begin
            addr_4_5 <= 13'h0;
          end else begin
            addr_4_5 <= (addr_4_5 + 13'h0001);
          end
        end
        if(weav_4_6) begin
          if(when_Weight_l326_70) begin
            addr_4_6 <= 13'h0;
          end else begin
            addr_4_6 <= (addr_4_6 + 13'h0001);
          end
        end
        if(weav_4_7) begin
          if(when_Weight_l326_71) begin
            addr_4_7 <= 13'h0;
          end else begin
            addr_4_7 <= (addr_4_7 + 13'h0001);
          end
        end
        if(weav_4_8) begin
          if(when_Weight_l326_72) begin
            addr_4_8 <= 13'h0;
          end else begin
            addr_4_8 <= (addr_4_8 + 13'h0001);
          end
        end
        if(weav_4_9) begin
          if(when_Weight_l326_73) begin
            addr_4_9 <= 13'h0;
          end else begin
            addr_4_9 <= (addr_4_9 + 13'h0001);
          end
        end
        if(weav_4_10) begin
          if(when_Weight_l326_74) begin
            addr_4_10 <= 13'h0;
          end else begin
            addr_4_10 <= (addr_4_10 + 13'h0001);
          end
        end
        if(weav_4_11) begin
          if(when_Weight_l326_75) begin
            addr_4_11 <= 13'h0;
          end else begin
            addr_4_11 <= (addr_4_11 + 13'h0001);
          end
        end
        if(weav_4_12) begin
          if(when_Weight_l326_76) begin
            addr_4_12 <= 13'h0;
          end else begin
            addr_4_12 <= (addr_4_12 + 13'h0001);
          end
        end
        if(weav_4_13) begin
          if(when_Weight_l326_77) begin
            addr_4_13 <= 13'h0;
          end else begin
            addr_4_13 <= (addr_4_13 + 13'h0001);
          end
        end
        if(weav_4_14) begin
          if(when_Weight_l326_78) begin
            addr_4_14 <= 13'h0;
          end else begin
            addr_4_14 <= (addr_4_14 + 13'h0001);
          end
        end
        if(weav_4_15) begin
          if(when_Weight_l326_79) begin
            addr_4_15 <= 13'h0;
          end else begin
            addr_4_15 <= (addr_4_15 + 13'h0001);
          end
        end
        if(weav_5_0) begin
          if(when_Weight_l326_80) begin
            addr_5_0 <= 13'h0;
          end else begin
            addr_5_0 <= (addr_5_0 + 13'h0001);
          end
        end
        if(weav_5_1) begin
          if(when_Weight_l326_81) begin
            addr_5_1 <= 13'h0;
          end else begin
            addr_5_1 <= (addr_5_1 + 13'h0001);
          end
        end
        if(weav_5_2) begin
          if(when_Weight_l326_82) begin
            addr_5_2 <= 13'h0;
          end else begin
            addr_5_2 <= (addr_5_2 + 13'h0001);
          end
        end
        if(weav_5_3) begin
          if(when_Weight_l326_83) begin
            addr_5_3 <= 13'h0;
          end else begin
            addr_5_3 <= (addr_5_3 + 13'h0001);
          end
        end
        if(weav_5_4) begin
          if(when_Weight_l326_84) begin
            addr_5_4 <= 13'h0;
          end else begin
            addr_5_4 <= (addr_5_4 + 13'h0001);
          end
        end
        if(weav_5_5) begin
          if(when_Weight_l326_85) begin
            addr_5_5 <= 13'h0;
          end else begin
            addr_5_5 <= (addr_5_5 + 13'h0001);
          end
        end
        if(weav_5_6) begin
          if(when_Weight_l326_86) begin
            addr_5_6 <= 13'h0;
          end else begin
            addr_5_6 <= (addr_5_6 + 13'h0001);
          end
        end
        if(weav_5_7) begin
          if(when_Weight_l326_87) begin
            addr_5_7 <= 13'h0;
          end else begin
            addr_5_7 <= (addr_5_7 + 13'h0001);
          end
        end
        if(weav_5_8) begin
          if(when_Weight_l326_88) begin
            addr_5_8 <= 13'h0;
          end else begin
            addr_5_8 <= (addr_5_8 + 13'h0001);
          end
        end
        if(weav_5_9) begin
          if(when_Weight_l326_89) begin
            addr_5_9 <= 13'h0;
          end else begin
            addr_5_9 <= (addr_5_9 + 13'h0001);
          end
        end
        if(weav_5_10) begin
          if(when_Weight_l326_90) begin
            addr_5_10 <= 13'h0;
          end else begin
            addr_5_10 <= (addr_5_10 + 13'h0001);
          end
        end
        if(weav_5_11) begin
          if(when_Weight_l326_91) begin
            addr_5_11 <= 13'h0;
          end else begin
            addr_5_11 <= (addr_5_11 + 13'h0001);
          end
        end
        if(weav_5_12) begin
          if(when_Weight_l326_92) begin
            addr_5_12 <= 13'h0;
          end else begin
            addr_5_12 <= (addr_5_12 + 13'h0001);
          end
        end
        if(weav_5_13) begin
          if(when_Weight_l326_93) begin
            addr_5_13 <= 13'h0;
          end else begin
            addr_5_13 <= (addr_5_13 + 13'h0001);
          end
        end
        if(weav_5_14) begin
          if(when_Weight_l326_94) begin
            addr_5_14 <= 13'h0;
          end else begin
            addr_5_14 <= (addr_5_14 + 13'h0001);
          end
        end
        if(weav_5_15) begin
          if(when_Weight_l326_95) begin
            addr_5_15 <= 13'h0;
          end else begin
            addr_5_15 <= (addr_5_15 + 13'h0001);
          end
        end
        if(weav_6_0) begin
          if(when_Weight_l326_96) begin
            addr_6_0 <= 13'h0;
          end else begin
            addr_6_0 <= (addr_6_0 + 13'h0001);
          end
        end
        if(weav_6_1) begin
          if(when_Weight_l326_97) begin
            addr_6_1 <= 13'h0;
          end else begin
            addr_6_1 <= (addr_6_1 + 13'h0001);
          end
        end
        if(weav_6_2) begin
          if(when_Weight_l326_98) begin
            addr_6_2 <= 13'h0;
          end else begin
            addr_6_2 <= (addr_6_2 + 13'h0001);
          end
        end
        if(weav_6_3) begin
          if(when_Weight_l326_99) begin
            addr_6_3 <= 13'h0;
          end else begin
            addr_6_3 <= (addr_6_3 + 13'h0001);
          end
        end
        if(weav_6_4) begin
          if(when_Weight_l326_100) begin
            addr_6_4 <= 13'h0;
          end else begin
            addr_6_4 <= (addr_6_4 + 13'h0001);
          end
        end
        if(weav_6_5) begin
          if(when_Weight_l326_101) begin
            addr_6_5 <= 13'h0;
          end else begin
            addr_6_5 <= (addr_6_5 + 13'h0001);
          end
        end
        if(weav_6_6) begin
          if(when_Weight_l326_102) begin
            addr_6_6 <= 13'h0;
          end else begin
            addr_6_6 <= (addr_6_6 + 13'h0001);
          end
        end
        if(weav_6_7) begin
          if(when_Weight_l326_103) begin
            addr_6_7 <= 13'h0;
          end else begin
            addr_6_7 <= (addr_6_7 + 13'h0001);
          end
        end
        if(weav_6_8) begin
          if(when_Weight_l326_104) begin
            addr_6_8 <= 13'h0;
          end else begin
            addr_6_8 <= (addr_6_8 + 13'h0001);
          end
        end
        if(weav_6_9) begin
          if(when_Weight_l326_105) begin
            addr_6_9 <= 13'h0;
          end else begin
            addr_6_9 <= (addr_6_9 + 13'h0001);
          end
        end
        if(weav_6_10) begin
          if(when_Weight_l326_106) begin
            addr_6_10 <= 13'h0;
          end else begin
            addr_6_10 <= (addr_6_10 + 13'h0001);
          end
        end
        if(weav_6_11) begin
          if(when_Weight_l326_107) begin
            addr_6_11 <= 13'h0;
          end else begin
            addr_6_11 <= (addr_6_11 + 13'h0001);
          end
        end
        if(weav_6_12) begin
          if(when_Weight_l326_108) begin
            addr_6_12 <= 13'h0;
          end else begin
            addr_6_12 <= (addr_6_12 + 13'h0001);
          end
        end
        if(weav_6_13) begin
          if(when_Weight_l326_109) begin
            addr_6_13 <= 13'h0;
          end else begin
            addr_6_13 <= (addr_6_13 + 13'h0001);
          end
        end
        if(weav_6_14) begin
          if(when_Weight_l326_110) begin
            addr_6_14 <= 13'h0;
          end else begin
            addr_6_14 <= (addr_6_14 + 13'h0001);
          end
        end
        if(weav_6_15) begin
          if(when_Weight_l326_111) begin
            addr_6_15 <= 13'h0;
          end else begin
            addr_6_15 <= (addr_6_15 + 13'h0001);
          end
        end
        if(weav_7_0) begin
          if(when_Weight_l326_112) begin
            addr_7_0 <= 13'h0;
          end else begin
            addr_7_0 <= (addr_7_0 + 13'h0001);
          end
        end
        if(weav_7_1) begin
          if(when_Weight_l326_113) begin
            addr_7_1 <= 13'h0;
          end else begin
            addr_7_1 <= (addr_7_1 + 13'h0001);
          end
        end
        if(weav_7_2) begin
          if(when_Weight_l326_114) begin
            addr_7_2 <= 13'h0;
          end else begin
            addr_7_2 <= (addr_7_2 + 13'h0001);
          end
        end
        if(weav_7_3) begin
          if(when_Weight_l326_115) begin
            addr_7_3 <= 13'h0;
          end else begin
            addr_7_3 <= (addr_7_3 + 13'h0001);
          end
        end
        if(weav_7_4) begin
          if(when_Weight_l326_116) begin
            addr_7_4 <= 13'h0;
          end else begin
            addr_7_4 <= (addr_7_4 + 13'h0001);
          end
        end
        if(weav_7_5) begin
          if(when_Weight_l326_117) begin
            addr_7_5 <= 13'h0;
          end else begin
            addr_7_5 <= (addr_7_5 + 13'h0001);
          end
        end
        if(weav_7_6) begin
          if(when_Weight_l326_118) begin
            addr_7_6 <= 13'h0;
          end else begin
            addr_7_6 <= (addr_7_6 + 13'h0001);
          end
        end
        if(weav_7_7) begin
          if(when_Weight_l326_119) begin
            addr_7_7 <= 13'h0;
          end else begin
            addr_7_7 <= (addr_7_7 + 13'h0001);
          end
        end
        if(weav_7_8) begin
          if(when_Weight_l326_120) begin
            addr_7_8 <= 13'h0;
          end else begin
            addr_7_8 <= (addr_7_8 + 13'h0001);
          end
        end
        if(weav_7_9) begin
          if(when_Weight_l326_121) begin
            addr_7_9 <= 13'h0;
          end else begin
            addr_7_9 <= (addr_7_9 + 13'h0001);
          end
        end
        if(weav_7_10) begin
          if(when_Weight_l326_122) begin
            addr_7_10 <= 13'h0;
          end else begin
            addr_7_10 <= (addr_7_10 + 13'h0001);
          end
        end
        if(weav_7_11) begin
          if(when_Weight_l326_123) begin
            addr_7_11 <= 13'h0;
          end else begin
            addr_7_11 <= (addr_7_11 + 13'h0001);
          end
        end
        if(weav_7_12) begin
          if(when_Weight_l326_124) begin
            addr_7_12 <= 13'h0;
          end else begin
            addr_7_12 <= (addr_7_12 + 13'h0001);
          end
        end
        if(weav_7_13) begin
          if(when_Weight_l326_125) begin
            addr_7_13 <= 13'h0;
          end else begin
            addr_7_13 <= (addr_7_13 + 13'h0001);
          end
        end
        if(weav_7_14) begin
          if(when_Weight_l326_126) begin
            addr_7_14 <= 13'h0;
          end else begin
            addr_7_14 <= (addr_7_14 + 13'h0001);
          end
        end
        if(weav_7_15) begin
          if(when_Weight_l326_127) begin
            addr_7_15 <= 13'h0;
          end else begin
            addr_7_15 <= (addr_7_15 + 13'h0001);
          end
        end
        if(weav_8_0) begin
          if(when_Weight_l326_128) begin
            addr_8_0 <= 13'h0;
          end else begin
            addr_8_0 <= (addr_8_0 + 13'h0001);
          end
        end
        if(weav_8_1) begin
          if(when_Weight_l326_129) begin
            addr_8_1 <= 13'h0;
          end else begin
            addr_8_1 <= (addr_8_1 + 13'h0001);
          end
        end
        if(weav_8_2) begin
          if(when_Weight_l326_130) begin
            addr_8_2 <= 13'h0;
          end else begin
            addr_8_2 <= (addr_8_2 + 13'h0001);
          end
        end
        if(weav_8_3) begin
          if(when_Weight_l326_131) begin
            addr_8_3 <= 13'h0;
          end else begin
            addr_8_3 <= (addr_8_3 + 13'h0001);
          end
        end
        if(weav_8_4) begin
          if(when_Weight_l326_132) begin
            addr_8_4 <= 13'h0;
          end else begin
            addr_8_4 <= (addr_8_4 + 13'h0001);
          end
        end
        if(weav_8_5) begin
          if(when_Weight_l326_133) begin
            addr_8_5 <= 13'h0;
          end else begin
            addr_8_5 <= (addr_8_5 + 13'h0001);
          end
        end
        if(weav_8_6) begin
          if(when_Weight_l326_134) begin
            addr_8_6 <= 13'h0;
          end else begin
            addr_8_6 <= (addr_8_6 + 13'h0001);
          end
        end
        if(weav_8_7) begin
          if(when_Weight_l326_135) begin
            addr_8_7 <= 13'h0;
          end else begin
            addr_8_7 <= (addr_8_7 + 13'h0001);
          end
        end
        if(weav_8_8) begin
          if(when_Weight_l326_136) begin
            addr_8_8 <= 13'h0;
          end else begin
            addr_8_8 <= (addr_8_8 + 13'h0001);
          end
        end
        if(weav_8_9) begin
          if(when_Weight_l326_137) begin
            addr_8_9 <= 13'h0;
          end else begin
            addr_8_9 <= (addr_8_9 + 13'h0001);
          end
        end
        if(weav_8_10) begin
          if(when_Weight_l326_138) begin
            addr_8_10 <= 13'h0;
          end else begin
            addr_8_10 <= (addr_8_10 + 13'h0001);
          end
        end
        if(weav_8_11) begin
          if(when_Weight_l326_139) begin
            addr_8_11 <= 13'h0;
          end else begin
            addr_8_11 <= (addr_8_11 + 13'h0001);
          end
        end
        if(weav_8_12) begin
          if(when_Weight_l326_140) begin
            addr_8_12 <= 13'h0;
          end else begin
            addr_8_12 <= (addr_8_12 + 13'h0001);
          end
        end
        if(weav_8_13) begin
          if(when_Weight_l326_141) begin
            addr_8_13 <= 13'h0;
          end else begin
            addr_8_13 <= (addr_8_13 + 13'h0001);
          end
        end
        if(weav_8_14) begin
          if(when_Weight_l326_142) begin
            addr_8_14 <= 13'h0;
          end else begin
            addr_8_14 <= (addr_8_14 + 13'h0001);
          end
        end
        if(weav_8_15) begin
          if(when_Weight_l326_143) begin
            addr_8_15 <= 13'h0;
          end else begin
            addr_8_15 <= (addr_8_15 + 13'h0001);
          end
        end
        if(when_WaCounter_l17_4) begin
          copyBias_copyCnt_count <= (copyBias_copyCnt_count + 8'h01);
          if(copyBias_copyCnt_valid) begin
            copyBias_copyCnt_count <= 8'h0;
          end
        end
        if(when_WaCounter_l17_5) begin
          copyScale_copyCnt_count <= (copyScale_copyCnt_count + 8'h01);
          if(copyScale_copyCnt_valid) begin
            copyScale_copyCnt_count <= 8'h0;
          end
        end
        if(when_WaCounter_l17_6) begin
          copyShift_copyCnt_count <= (copyShift_copyCnt_count + 8'h01);
          if(copyShift_copyCnt_valid) begin
            copyShift_copyCnt_count <= 8'h0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    channelInTimes <= (channelIn >>> 4);
    channelOutTimes <= channelOut;
    case(convType)
      2'b10 : begin
        copyTimes <= 4'b0000;
      end
      2'b01 : begin
        copyTimes <= 4'b0111;
      end
      default : begin
        copyTimes <= 4'b0000;
      end
    endcase
  end


endmodule

module ConvComputeCtrl (
  input               start,
  output reg          mDataValid,
  input               mDataReady,
  output              normPreValid,
  input               sDataReady,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input      [11:0]   channelIn,
  input      [11:0]   channelOut,
  output     [4:0]    featureMemReadAddr,
  output     [4:0]    featureMemWriteAddr,
  output reg          featureMemWriteReady,
  output     [8:0]    weightReadAddr_0,
  output     [8:0]    weightReadAddr_1,
  output     [8:0]    weightReadAddr_2,
  output     [8:0]    weightReadAddr_3,
  output     [8:0]    weightReadAddr_4,
  output     [8:0]    weightReadAddr_5,
  output     [8:0]    weightReadAddr_6,
  output     [8:0]    weightReadAddr_7,
  output     [8:0]    weightReadAddr_8,
  output     [5:0]    biasReadAddr,
  output     [5:0]    scaleReadAddr,
  output     [5:0]    shiftReadAddr,
  input               activationEn,
  output     [12:0]   sCount,
  output     [12:0]   mCount,
  input      [1:0]    convType,
  input               clk,
  input               reset,
  input               softReset
);
  localparam ConvComputeCtrlEnum_IDLE = 6'd1;
  localparam ConvComputeCtrlEnum_INIT = 6'd2;
  localparam ConvComputeCtrlEnum_DATA_READY = 6'd4;
  localparam ConvComputeCtrlEnum_FIFO_READY = 6'd8;
  localparam ConvComputeCtrlEnum_COMPUTE = 6'd16;
  localparam ConvComputeCtrlEnum_END_1 = 6'd32;

  wire       [7:0]    _zz_temp;
  wire       [4:0]    _zz_temp_1;
  wire       [11:0]   _zz_when_WaCounter_l12_1;
  wire       [11:0]   _zz_when_WaCounter_l12_2;
  wire       [7:0]    _zz_when_WaCounter_l12_2_1;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire       [9:0]    _zz_when_WaCounter_l12_4;
  wire       [7:0]    _zz_when_WaCounter_l12_5;
  wire       [7:0]    _zz_when_WaCounter_l12_5_1;
  wire                convComputeCtrlFsm_start;
  wire                convComputeCtrlFsm_dataReady;
  wire                convComputeCtrlFsm_fifoReady;
  reg                 convComputeCtrlFsm_initEnd;
  reg                 convComputeCtrlFsm_computeEnd;
  reg                 convComputeCtrlFsm_endEnd;
  reg        [5:0]    convComputeCtrlFsm_currentState;
  reg        [5:0]    convComputeCtrlFsm_nextState;
  wire                when_WaCounter_l17;
  reg        [2:0]    initCnt_count;
  reg                 initCnt_valid;
  wire                when_WaCounter_l12;
  reg        [11:0]   temp;
  reg        [11:0]   channelInTimes;
  reg        [7:0]    channelOutTimes;
  wire                when_WaCounter_l17_1;
  reg        [11:0]   channelInCnt_count;
  reg                 channelInCnt_valid;
  wire                when_WaCounter_l12_1;
  wire                when_WaCounter_l17_2;
  reg        [11:0]   channelOutCnt_count;
  reg                 channelOutCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                when_WaCounter_l17_3;
  reg        [9:0]    columnCnt_count;
  reg                 columnCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                when_WaCounter_l17_4;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_4;
  wire                when_ConvComputeCtrl_l137;
  wire                when_WaUtil_l29;
  wire                when_WaUtil_l29_1;
  (* max_fanout = "50" *) reg        [4:0]    featureMemWriteAddr_1;
  wire                when_ConvComputeCtrl_l150;
  (* max_fanout = "50" *) reg        [4:0]    featureMemReadAddrTemp;
  wire                when_ConvComputeCtrl_l159;
  reg        [4:0]    featureMemReadAddrTemp_delay_1;
  (* max_fanout = "50" *) reg        [4:0]    featureMemReadAddrTemp_delay_2;
  (* max_fanout = "50" *) reg        [8:0]    weightReadAddr;
  wire                when_ConvComputeCtrl_l160;
  wire                when_ConvComputeCtrl_l159_1;
  (* max_fanout = "50" *) reg        [8:0]    weightReadAddrTemp;
  reg                 channelTimesAdd;
  wire                when_WaUtil_l29_2;
  reg                 channelTimesAdd_delay_1;
  reg                 channelTimesAdd_delay_2;
  reg                 channelTimesAdd_delay_3;
  reg                 channelTimesAdd_delay_4;
  reg                 channelTimesAdd_delay_5;
  reg                 channelTimesAdd_delay_6;
  reg                 channelTimesAdd_delay_7;
  reg                 channelTimesAdd_delay_8;
  reg                 channelTimesAdd_delay_9;
  reg                 channelTimesAdd_delay_10;
  reg                 channelTimesAdd_delay_11;
  reg                 channelTimesAdd_delay_12;
  reg                 channelTimesAdd_delay_13;
  reg                 channelTimesAdd_delay_14;
  reg                 channelTimesAdd_delay_15;
  reg                 channelTimesAdd_delay_16;
  reg                 channelTimesAdd_delay_17;
  reg                 channelTimesAdd_delay_18;
  reg                 channelTimesAdd_delay_19;
  reg                 channelTimesAdd_delay_20;
  reg                 channelTimesAdd_delay_21;
  reg                 channelTimesAdd_delay_22;
  reg                 channelTimesAdd_delay_23;
  reg                 channelTimesAdd_delay_24;
  reg                 channelTimesAdd_delay_25;
  reg                 channelTimesAdd_delay_26;
  reg                 normValidTemp;
  wire                when_WaUtil_l29_3;
  wire                normValidTempQ_0;
  reg                 normValidTempQ_1;
  reg                 normValidTempQ_2;
  reg                 normValidTempQ_3;
  reg                 normValidTempQ_4;
  reg                 normValidTempQ_5;
  reg                 normValidTempQ_6;
  reg                 normValidTempQ_7;
  reg                 normValidTempQ_8;
  reg                 normValidTempQ_9;
  reg                 normValidTempQ_10;
  reg                 normValidTempQ_11;
  reg                 normValidTempQ_12;
  reg                 normValidTempQ_13;
  reg                 normValidTempQ_14;
  reg                 normValidTempQ_15;
  reg                 normValidTempQ_16;
  reg                 normValidTempQ_17;
  reg                 normValidTempQ_18;
  reg                 normValidTempQ_19;
  reg                 normValidTempQ_20;
  reg                 normValidTempQ_21;
  reg                 normValidTempQ_22;
  reg                 normValidTempQ_23;
  reg                 normValidTempQ_24;
  reg                 normValidTempQ_25;
  reg                 normValidTempQ_26;
  reg                 normValidTempQ_27;
  reg                 normValidTempQ_28;
  reg                 normValidTempQ_29;
  reg                 normValidTempQ_30;
  reg                 normValidTempQ_31;
  reg                 normValidTempQ_32;
  reg                 normValidTempQ_33;
  reg                 normValidTempQ_34;
  reg                 normValidTempQ_35;
  reg                 normValidTempQ_36;
  reg                 normValidTempQ_37;
  reg                 normValidTempQ_38;
  reg                 normValidTempQ_39;
  reg                 normValidTempQ_40;
  reg                 normValidTempQ_41;
  reg                 normValidTempQ_42;
  reg                 normValidTempQ_43;
  reg                 normValidTempQ_44;
  reg                 normValidTempQ_45;
  reg                 normValidTempQ_46;
  reg                 normValidTempQ_47;
  reg                 normValidTempQ_48;
  reg                 normValidTempQ_49;
  reg                 normValidTempQ_50;
  reg        [21:0]   _zz_sCount;
  reg        [5:0]    biasAddrCnt_count;
  reg                 biasAddrCnt_valid;
  wire                when_WaCounter_l12_5;
  `ifndef SYNTHESIS
  reg [79:0] convComputeCtrlFsm_currentState_string;
  reg [79:0] convComputeCtrlFsm_nextState_string;
  `endif


  assign _zz_temp = (channelIn >>> 4);
  assign _zz_temp_1 = (channelIn >>> 7);
  assign _zz_when_WaCounter_l12_1 = (channelInTimes - 12'h001);
  assign _zz_when_WaCounter_l12_2_1 = (channelOutTimes - 8'h01);
  assign _zz_when_WaCounter_l12_2 = {4'd0, _zz_when_WaCounter_l12_2_1};
  assign _zz_when_WaCounter_l12_3 = (colNumIn - 10'h001);
  assign _zz_when_WaCounter_l12_4 = (rowNumIn - 10'h001);
  assign _zz_when_WaCounter_l12_5 = {2'd0, biasAddrCnt_count};
  assign _zz_when_WaCounter_l12_5_1 = (channelOutTimes - 8'h01);
  `ifndef SYNTHESIS
  always @(*) begin
    case(convComputeCtrlFsm_currentState)
      ConvComputeCtrlEnum_IDLE : convComputeCtrlFsm_currentState_string = "IDLE      ";
      ConvComputeCtrlEnum_INIT : convComputeCtrlFsm_currentState_string = "INIT      ";
      ConvComputeCtrlEnum_DATA_READY : convComputeCtrlFsm_currentState_string = "DATA_READY";
      ConvComputeCtrlEnum_FIFO_READY : convComputeCtrlFsm_currentState_string = "FIFO_READY";
      ConvComputeCtrlEnum_COMPUTE : convComputeCtrlFsm_currentState_string = "COMPUTE   ";
      ConvComputeCtrlEnum_END_1 : convComputeCtrlFsm_currentState_string = "END_1     ";
      default : convComputeCtrlFsm_currentState_string = "??????????";
    endcase
  end
  always @(*) begin
    case(convComputeCtrlFsm_nextState)
      ConvComputeCtrlEnum_IDLE : convComputeCtrlFsm_nextState_string = "IDLE      ";
      ConvComputeCtrlEnum_INIT : convComputeCtrlFsm_nextState_string = "INIT      ";
      ConvComputeCtrlEnum_DATA_READY : convComputeCtrlFsm_nextState_string = "DATA_READY";
      ConvComputeCtrlEnum_FIFO_READY : convComputeCtrlFsm_nextState_string = "FIFO_READY";
      ConvComputeCtrlEnum_COMPUTE : convComputeCtrlFsm_nextState_string = "COMPUTE   ";
      ConvComputeCtrlEnum_END_1 : convComputeCtrlFsm_nextState_string = "END_1     ";
      default : convComputeCtrlFsm_nextState_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((convComputeCtrlFsm_currentState) & ConvComputeCtrlEnum_IDLE) == ConvComputeCtrlEnum_IDLE) : begin
        if(convComputeCtrlFsm_start) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_INIT;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_IDLE;
        end
      end
      (((convComputeCtrlFsm_currentState) & ConvComputeCtrlEnum_INIT) == ConvComputeCtrlEnum_INIT) : begin
        if(convComputeCtrlFsm_initEnd) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_DATA_READY;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_INIT;
        end
      end
      (((convComputeCtrlFsm_currentState) & ConvComputeCtrlEnum_DATA_READY) == ConvComputeCtrlEnum_DATA_READY) : begin
        if(convComputeCtrlFsm_dataReady) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_FIFO_READY;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_DATA_READY;
        end
      end
      (((convComputeCtrlFsm_currentState) & ConvComputeCtrlEnum_FIFO_READY) == ConvComputeCtrlEnum_FIFO_READY) : begin
        if(convComputeCtrlFsm_fifoReady) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_COMPUTE;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_FIFO_READY;
        end
      end
      (((convComputeCtrlFsm_currentState) & ConvComputeCtrlEnum_COMPUTE) == ConvComputeCtrlEnum_COMPUTE) : begin
        if(convComputeCtrlFsm_computeEnd) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_END_1;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_COMPUTE;
        end
      end
      default : begin
        if(convComputeCtrlFsm_endEnd) begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_IDLE;
        end else begin
          convComputeCtrlFsm_nextState = ConvComputeCtrlEnum_DATA_READY;
        end
      end
    endcase
  end

  assign convComputeCtrlFsm_start = start;
  assign convComputeCtrlFsm_dataReady = sDataReady;
  assign convComputeCtrlFsm_fifoReady = mDataReady;
  assign when_WaCounter_l17 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_INIT) != 6'b000000);
  assign when_WaCounter_l12 = (initCnt_count == 3'b111);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCnt_valid = 1'b1;
    end else begin
      initCnt_valid = 1'b0;
    end
  end

  always @(*) begin
    case(convType)
      2'b00, 2'b10 : begin
        temp = {4'd0, _zz_temp};
      end
      2'b01 : begin
        temp = {7'd0, _zz_temp_1};
      end
      default : begin
        temp = 12'h0;
      end
    endcase
  end

  assign when_WaCounter_l17_1 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000);
  assign when_WaCounter_l12_1 = (channelInCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelInCnt_valid = 1'b1;
    end else begin
      channelInCnt_valid = 1'b0;
    end
    if(when_ConvComputeCtrl_l137) begin
      channelInCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_2 = (((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000) && channelInCnt_valid);
  assign when_WaCounter_l12_2 = (channelOutCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      channelOutCnt_valid = 1'b1;
    end else begin
      channelOutCnt_valid = 1'b0;
    end
    if(when_ConvComputeCtrl_l137) begin
      channelOutCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_3 = ((((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000) && channelInCnt_valid) && channelOutCnt_valid);
  assign when_WaCounter_l12_3 = (columnCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      columnCnt_valid = 1'b1;
    end else begin
      columnCnt_valid = 1'b0;
    end
    if(when_ConvComputeCtrl_l137) begin
      columnCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_4 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_END_1) != 6'b000000);
  assign when_WaCounter_l12_4 = (rowCnt_count == _zz_when_WaCounter_l12_4);
  always @(*) begin
    if(when_WaCounter_l12_4) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
  end

  assign when_ConvComputeCtrl_l137 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_IDLE) != 6'b000000);
  assign when_WaUtil_l29 = ((channelInCnt_valid && channelOutCnt_valid) && columnCnt_valid);
  always @(*) begin
    if(when_WaUtil_l29) begin
      convComputeCtrlFsm_computeEnd = 1'b1;
    end else begin
      convComputeCtrlFsm_computeEnd = 1'b0;
    end
  end

  always @(*) begin
    if(rowCnt_valid) begin
      convComputeCtrlFsm_endEnd = 1'b1;
    end else begin
      convComputeCtrlFsm_endEnd = 1'b0;
    end
  end

  always @(*) begin
    if(initCnt_valid) begin
      convComputeCtrlFsm_initEnd = 1'b1;
    end else begin
      convComputeCtrlFsm_initEnd = 1'b0;
    end
  end

  assign when_WaUtil_l29_1 = (((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000) && (channelOutCnt_count == 12'h0));
  assign featureMemWriteAddr = featureMemWriteAddr_1;
  assign when_ConvComputeCtrl_l150 = ((channelOutCnt_count == 12'h0) && (channelInCnt_count == 12'h0));
  assign when_ConvComputeCtrl_l159 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000);
  assign featureMemReadAddr = featureMemReadAddrTemp_delay_2;
  assign when_ConvComputeCtrl_l160 = (channelInCnt_valid && channelOutCnt_valid);
  assign when_ConvComputeCtrl_l159_1 = ((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000);
  assign weightReadAddr_0 = weightReadAddrTemp;
  assign weightReadAddr_1 = weightReadAddrTemp;
  assign weightReadAddr_2 = weightReadAddrTemp;
  assign weightReadAddr_3 = weightReadAddrTemp;
  assign weightReadAddr_4 = weightReadAddrTemp;
  assign weightReadAddr_5 = weightReadAddrTemp;
  assign weightReadAddr_6 = weightReadAddrTemp;
  assign weightReadAddr_7 = weightReadAddrTemp;
  assign weightReadAddr_8 = weightReadAddrTemp;
  assign when_WaUtil_l29_2 = (((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000) && (channelInCnt_count == 12'h0));
  assign normPreValid = channelTimesAdd_delay_26;
  assign when_WaUtil_l29_3 = (((convComputeCtrlFsm_currentState & ConvComputeCtrlEnum_COMPUTE) != 6'b000000) && channelInCnt_valid);
  assign normValidTempQ_0 = normValidTemp;
  assign sCount = _zz_sCount[12:0];
  assign mCount = sCount;
  assign when_WaCounter_l12_5 = (_zz_when_WaCounter_l12_5 == _zz_when_WaCounter_l12_5_1);
  always @(*) begin
    if(when_WaCounter_l12_5) begin
      biasAddrCnt_valid = 1'b1;
    end else begin
      biasAddrCnt_valid = 1'b0;
    end
  end

  assign biasReadAddr = biasAddrCnt_count;
  assign scaleReadAddr = biasAddrCnt_count;
  assign shiftReadAddr = biasAddrCnt_count;
  always @(*) begin
    if(activationEn) begin
      mDataValid = normValidTempQ_50;
    end else begin
      mDataValid = normValidTempQ_42;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      featureMemWriteReady <= 1'b0;
      convComputeCtrlFsm_currentState <= ConvComputeCtrlEnum_IDLE;
      initCnt_count <= 3'b000;
      channelInCnt_count <= 12'h0;
      channelOutCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      featureMemWriteAddr_1 <= 5'h0;
      featureMemReadAddrTemp <= 5'h0;
      channelTimesAdd <= 1'b0;
      normValidTemp <= 1'b0;
      biasAddrCnt_count <= 6'h0;
    end else begin
      if(softReset) begin
      featureMemWriteReady <= 1'b0;
      convComputeCtrlFsm_currentState <= ConvComputeCtrlEnum_IDLE;
      initCnt_count <= 3'b000;
      channelInCnt_count <= 12'h0;
      channelOutCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      featureMemWriteAddr_1 <= 5'h0;
      featureMemReadAddrTemp <= 5'h0;
      channelTimesAdd <= 1'b0;
      normValidTemp <= 1'b0;
      biasAddrCnt_count <= 6'h0;
      end else begin
        convComputeCtrlFsm_currentState <= convComputeCtrlFsm_nextState;
        if(when_WaCounter_l17) begin
          initCnt_count <= (initCnt_count + 3'b001);
          if(initCnt_valid) begin
            initCnt_count <= 3'b000;
          end
        end
        if(when_WaCounter_l17_1) begin
          channelInCnt_count <= (channelInCnt_count + 12'h001);
          if(channelInCnt_valid) begin
            channelInCnt_count <= 12'h0;
          end
        end
        if(when_WaCounter_l17_2) begin
          channelOutCnt_count <= (channelOutCnt_count + 12'h001);
          if(channelOutCnt_valid) begin
            channelOutCnt_count <= 12'h0;
          end
        end
        if(when_WaCounter_l17_3) begin
          columnCnt_count <= (columnCnt_count + 10'h001);
          if(columnCnt_valid) begin
            columnCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_4) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
        if(when_ConvComputeCtrl_l137) begin
          channelInCnt_count <= 12'h0;
          channelOutCnt_count <= 12'h0;
          columnCnt_count <= 10'h0;
        end
        if(when_WaUtil_l29_1) begin
          featureMemWriteReady <= 1'b1;
        end else begin
          featureMemWriteReady <= 1'b0;
        end
        if(when_ConvComputeCtrl_l150) begin
          featureMemWriteAddr_1 <= 5'h0;
        end else begin
          if(featureMemWriteReady) begin
            featureMemWriteAddr_1 <= (featureMemWriteAddr_1 + 5'h01);
          end else begin
            featureMemWriteAddr_1 <= 5'h0;
          end
        end
        if(when_ConvComputeCtrl_l159) begin
          if(channelInCnt_valid) begin
            featureMemReadAddrTemp <= 5'h0;
          end else begin
            featureMemReadAddrTemp <= (featureMemReadAddrTemp + 5'h01);
          end
        end else begin
          featureMemReadAddrTemp <= 5'h0;
        end
        if(when_WaUtil_l29_2) begin
          channelTimesAdd <= 1'b1;
        end else begin
          channelTimesAdd <= 1'b0;
        end
        if(when_WaUtil_l29_3) begin
          normValidTemp <= 1'b1;
        end else begin
          normValidTemp <= 1'b0;
        end
        if(normValidTempQ_26) begin
          biasAddrCnt_count <= (biasAddrCnt_count + 6'h01);
          if(biasAddrCnt_valid) begin
            biasAddrCnt_count <= 6'h0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    channelInTimes <= temp;
    channelOutTimes <= (channelOut >>> 4);
    featureMemReadAddrTemp_delay_1 <= featureMemReadAddrTemp;
    featureMemReadAddrTemp_delay_2 <= featureMemReadAddrTemp_delay_1;
    if(when_ConvComputeCtrl_l159_1) begin
      if(when_ConvComputeCtrl_l160) begin
        weightReadAddr <= 9'h0;
      end else begin
        weightReadAddr <= (weightReadAddr + 9'h001);
      end
    end else begin
      weightReadAddr <= 9'h0;
    end
    weightReadAddrTemp <= weightReadAddr;
    channelTimesAdd_delay_1 <= channelTimesAdd;
    channelTimesAdd_delay_2 <= channelTimesAdd_delay_1;
    channelTimesAdd_delay_3 <= channelTimesAdd_delay_2;
    channelTimesAdd_delay_4 <= channelTimesAdd_delay_3;
    channelTimesAdd_delay_5 <= channelTimesAdd_delay_4;
    channelTimesAdd_delay_6 <= channelTimesAdd_delay_5;
    channelTimesAdd_delay_7 <= channelTimesAdd_delay_6;
    channelTimesAdd_delay_8 <= channelTimesAdd_delay_7;
    channelTimesAdd_delay_9 <= channelTimesAdd_delay_8;
    channelTimesAdd_delay_10 <= channelTimesAdd_delay_9;
    channelTimesAdd_delay_11 <= channelTimesAdd_delay_10;
    channelTimesAdd_delay_12 <= channelTimesAdd_delay_11;
    channelTimesAdd_delay_13 <= channelTimesAdd_delay_12;
    channelTimesAdd_delay_14 <= channelTimesAdd_delay_13;
    channelTimesAdd_delay_15 <= channelTimesAdd_delay_14;
    channelTimesAdd_delay_16 <= channelTimesAdd_delay_15;
    channelTimesAdd_delay_17 <= channelTimesAdd_delay_16;
    channelTimesAdd_delay_18 <= channelTimesAdd_delay_17;
    channelTimesAdd_delay_19 <= channelTimesAdd_delay_18;
    channelTimesAdd_delay_20 <= channelTimesAdd_delay_19;
    channelTimesAdd_delay_21 <= channelTimesAdd_delay_20;
    channelTimesAdd_delay_22 <= channelTimesAdd_delay_21;
    channelTimesAdd_delay_23 <= channelTimesAdd_delay_22;
    channelTimesAdd_delay_24 <= channelTimesAdd_delay_23;
    channelTimesAdd_delay_25 <= channelTimesAdd_delay_24;
    channelTimesAdd_delay_26 <= channelTimesAdd_delay_25;
    normValidTempQ_1 <= normValidTempQ_0;
    normValidTempQ_2 <= normValidTempQ_1;
    normValidTempQ_3 <= normValidTempQ_2;
    normValidTempQ_4 <= normValidTempQ_3;
    normValidTempQ_5 <= normValidTempQ_4;
    normValidTempQ_6 <= normValidTempQ_5;
    normValidTempQ_7 <= normValidTempQ_6;
    normValidTempQ_8 <= normValidTempQ_7;
    normValidTempQ_9 <= normValidTempQ_8;
    normValidTempQ_10 <= normValidTempQ_9;
    normValidTempQ_11 <= normValidTempQ_10;
    normValidTempQ_12 <= normValidTempQ_11;
    normValidTempQ_13 <= normValidTempQ_12;
    normValidTempQ_14 <= normValidTempQ_13;
    normValidTempQ_15 <= normValidTempQ_14;
    normValidTempQ_16 <= normValidTempQ_15;
    normValidTempQ_17 <= normValidTempQ_16;
    normValidTempQ_18 <= normValidTempQ_17;
    normValidTempQ_19 <= normValidTempQ_18;
    normValidTempQ_20 <= normValidTempQ_19;
    normValidTempQ_21 <= normValidTempQ_20;
    normValidTempQ_22 <= normValidTempQ_21;
    normValidTempQ_23 <= normValidTempQ_22;
    normValidTempQ_24 <= normValidTempQ_23;
    normValidTempQ_25 <= normValidTempQ_24;
    normValidTempQ_26 <= normValidTempQ_25;
    normValidTempQ_27 <= normValidTempQ_26;
    normValidTempQ_28 <= normValidTempQ_27;
    normValidTempQ_29 <= normValidTempQ_28;
    normValidTempQ_30 <= normValidTempQ_29;
    normValidTempQ_31 <= normValidTempQ_30;
    normValidTempQ_32 <= normValidTempQ_31;
    normValidTempQ_33 <= normValidTempQ_32;
    normValidTempQ_34 <= normValidTempQ_33;
    normValidTempQ_35 <= normValidTempQ_34;
    normValidTempQ_36 <= normValidTempQ_35;
    normValidTempQ_37 <= normValidTempQ_36;
    normValidTempQ_38 <= normValidTempQ_37;
    normValidTempQ_39 <= normValidTempQ_38;
    normValidTempQ_40 <= normValidTempQ_39;
    normValidTempQ_41 <= normValidTempQ_40;
    normValidTempQ_42 <= normValidTempQ_41;
    normValidTempQ_43 <= normValidTempQ_42;
    normValidTempQ_44 <= normValidTempQ_43;
    normValidTempQ_45 <= normValidTempQ_44;
    normValidTempQ_46 <= normValidTempQ_45;
    normValidTempQ_47 <= normValidTempQ_46;
    normValidTempQ_48 <= normValidTempQ_47;
    normValidTempQ_49 <= normValidTempQ_48;
    normValidTempQ_50 <= normValidTempQ_49;
    _zz_sCount <= (colNumIn * channelInTimes);
  end


endmodule

module DataGenerate (
  input               sData_valid,
  output reg          sData_ready,
  input      [127:0]  sData_payload,
  input               start,
  input               enPadding,
  input      [11:0]   channelIn,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input      [7:0]    zeroDara,
  input      [0:0]    zeroNum,
  output reg          mData_mData_0_valid,
  output reg [127:0]  mData_mData_0_payload,
  output reg          mData_mData_1_valid,
  output reg [127:0]  mData_mData_1_payload,
  output reg          mData_mData_2_valid,
  output reg [127:0]  mData_mData_2_payload,
  output reg          mData_mData_3_valid,
  output reg [127:0]  mData_mData_3_payload,
  output reg          mData_mData_4_valid,
  output reg [127:0]  mData_mData_4_payload,
  output reg          mData_mData_5_valid,
  output reg [127:0]  mData_mData_5_payload,
  output reg          mData_mData_6_valid,
  output reg [127:0]  mData_mData_6_payload,
  output reg          mData_mData_7_valid,
  output reg [127:0]  mData_mData_7_payload,
  output reg          mData_mData_8_valid,
  output reg [127:0]  mData_mData_8_payload,
  input               mData_ready,
  input      [1:0]    convType,
  input               reset,
  input               clk,
  input               softReset
);

  reg                 padding_1_sData_valid;
  reg        [127:0]  padding_1_sData_payload;
  reg                 padding_1_start;
  reg                 featureGenerate_1_mData_ready;
  reg                 featureWidthConvert_1_sData_valid;
  reg        [127:0]  featureWidthConvert_1_sData_payload;
  reg                 featureWidthConvert_1_mData_ready;
  reg                 featureWidthConvert_1_start;
  reg                 featureConv11Convert_1_io_sData_valid;
  reg        [127:0]  featureConv11Convert_1_io_sData_payload;
  reg                 featureConv11Convert_1_io_mData_ready;
  reg                 featureConv11Convert_1_io_start;
  wire                padding_1_sData_ready;
  wire                padding_1_mData_valid;
  wire       [127:0]  padding_1_mData_payload;
  wire       [9:0]    padding_1_rowNumOut;
  wire       [9:0]    padding_1_colNumOut;
  wire                featureGenerate_1_sData_ready;
  wire                featureGenerate_1_mData_mData_0_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_0_payload;
  wire                featureGenerate_1_mData_mData_1_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_1_payload;
  wire                featureGenerate_1_mData_mData_2_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_2_payload;
  wire                featureGenerate_1_mData_mData_3_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_3_payload;
  wire                featureGenerate_1_mData_mData_4_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_4_payload;
  wire                featureGenerate_1_mData_mData_5_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_5_payload;
  wire                featureGenerate_1_mData_mData_6_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_6_payload;
  wire                featureGenerate_1_mData_mData_7_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_7_payload;
  wire                featureGenerate_1_mData_mData_8_valid;
  wire       [127:0]  featureGenerate_1_mData_mData_8_payload;
  wire                featureWidthConvert_1_sData_ready;
  wire                featureWidthConvert_1_mData_mData_0_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_0_payload;
  wire                featureWidthConvert_1_mData_mData_1_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_1_payload;
  wire                featureWidthConvert_1_mData_mData_2_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_2_payload;
  wire                featureWidthConvert_1_mData_mData_3_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_3_payload;
  wire                featureWidthConvert_1_mData_mData_4_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_4_payload;
  wire                featureWidthConvert_1_mData_mData_5_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_5_payload;
  wire                featureWidthConvert_1_mData_mData_6_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_6_payload;
  wire                featureWidthConvert_1_mData_mData_7_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_7_payload;
  wire                featureWidthConvert_1_mData_mData_8_valid;
  wire       [127:0]  featureWidthConvert_1_mData_mData_8_payload;
  wire                featureConv11Convert_1_io_sData_ready;
  wire                featureConv11Convert_1_io_mData_mData_0_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_0_payload;
  wire                featureConv11Convert_1_io_mData_mData_1_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_1_payload;
  wire                featureConv11Convert_1_io_mData_mData_2_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_2_payload;
  wire                featureConv11Convert_1_io_mData_mData_3_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_3_payload;
  wire                featureConv11Convert_1_io_mData_mData_4_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_4_payload;
  wire                featureConv11Convert_1_io_mData_mData_5_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_5_payload;
  wire                featureConv11Convert_1_io_mData_mData_6_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_6_payload;
  wire                featureConv11Convert_1_io_mData_mData_7_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_7_payload;
  wire                featureConv11Convert_1_io_mData_mData_8_valid;
  wire       [127:0]  featureConv11Convert_1_io_mData_mData_8_payload;

  Padding padding_1 (
    .sData_valid   (padding_1_sData_valid         ), //i
    .sData_ready   (padding_1_sData_ready         ), //o
    .sData_payload (padding_1_sData_payload[127:0]), //i
    .mData_valid   (padding_1_mData_valid         ), //o
    .mData_ready   (featureGenerate_1_sData_ready ), //i
    .mData_payload (padding_1_mData_payload[127:0]), //o
    .enPadding     (enPadding                     ), //i
    .channelIn     (channelIn[11:0]               ), //i
    .start         (padding_1_start               ), //i
    .rowNumIn      (rowNumIn[9:0]                 ), //i
    .rowNumOut     (padding_1_rowNumOut[9:0]      ), //o
    .colNumIn      (colNumIn[9:0]                 ), //i
    .colNumOut     (padding_1_colNumOut[9:0]      ), //o
    .zeroDara      (zeroDara[7:0]                 ), //i
    .zeroNum       (zeroNum                       ), //i
    .clk           (clk                           ), //i
    .reset         (reset                         ), //i
    .softReset     (softReset                     )  //i
  );
  FeatureGenerate featureGenerate_1 (
    .sData_valid           (padding_1_mData_valid                         ), //i
    .sData_ready           (featureGenerate_1_sData_ready                 ), //o
    .sData_payload         (padding_1_mData_payload[127:0]                ), //i
    .mData_mData_0_valid   (featureGenerate_1_mData_mData_0_valid         ), //o
    .mData_mData_0_payload (featureGenerate_1_mData_mData_0_payload[127:0]), //o
    .mData_mData_1_valid   (featureGenerate_1_mData_mData_1_valid         ), //o
    .mData_mData_1_payload (featureGenerate_1_mData_mData_1_payload[127:0]), //o
    .mData_mData_2_valid   (featureGenerate_1_mData_mData_2_valid         ), //o
    .mData_mData_2_payload (featureGenerate_1_mData_mData_2_payload[127:0]), //o
    .mData_mData_3_valid   (featureGenerate_1_mData_mData_3_valid         ), //o
    .mData_mData_3_payload (featureGenerate_1_mData_mData_3_payload[127:0]), //o
    .mData_mData_4_valid   (featureGenerate_1_mData_mData_4_valid         ), //o
    .mData_mData_4_payload (featureGenerate_1_mData_mData_4_payload[127:0]), //o
    .mData_mData_5_valid   (featureGenerate_1_mData_mData_5_valid         ), //o
    .mData_mData_5_payload (featureGenerate_1_mData_mData_5_payload[127:0]), //o
    .mData_mData_6_valid   (featureGenerate_1_mData_mData_6_valid         ), //o
    .mData_mData_6_payload (featureGenerate_1_mData_mData_6_payload[127:0]), //o
    .mData_mData_7_valid   (featureGenerate_1_mData_mData_7_valid         ), //o
    .mData_mData_7_payload (featureGenerate_1_mData_mData_7_payload[127:0]), //o
    .mData_mData_8_valid   (featureGenerate_1_mData_mData_8_valid         ), //o
    .mData_mData_8_payload (featureGenerate_1_mData_mData_8_payload[127:0]), //o
    .mData_ready           (featureGenerate_1_mData_ready                 ), //i
    .rowNumIn              (padding_1_rowNumOut[9:0]                      ), //i
    .colNumIn              (padding_1_colNumOut[9:0]                      ), //i
    .start                 (padding_1_start                               ), //i
    .channelIn             (channelIn[11:0]                               ), //i
    .clk                   (clk                                           ), //i
    .reset                 (reset                                         ), //i
    .softReset             (softReset                                     )  //i
  );
  FeatureWidthConvert featureWidthConvert_1 (
    .sData_valid           (featureWidthConvert_1_sData_valid                 ), //i
    .sData_ready           (featureWidthConvert_1_sData_ready                 ), //o
    .sData_payload         (featureWidthConvert_1_sData_payload[127:0]        ), //i
    .mData_mData_0_valid   (featureWidthConvert_1_mData_mData_0_valid         ), //o
    .mData_mData_0_payload (featureWidthConvert_1_mData_mData_0_payload[127:0]), //o
    .mData_mData_1_valid   (featureWidthConvert_1_mData_mData_1_valid         ), //o
    .mData_mData_1_payload (featureWidthConvert_1_mData_mData_1_payload[127:0]), //o
    .mData_mData_2_valid   (featureWidthConvert_1_mData_mData_2_valid         ), //o
    .mData_mData_2_payload (featureWidthConvert_1_mData_mData_2_payload[127:0]), //o
    .mData_mData_3_valid   (featureWidthConvert_1_mData_mData_3_valid         ), //o
    .mData_mData_3_payload (featureWidthConvert_1_mData_mData_3_payload[127:0]), //o
    .mData_mData_4_valid   (featureWidthConvert_1_mData_mData_4_valid         ), //o
    .mData_mData_4_payload (featureWidthConvert_1_mData_mData_4_payload[127:0]), //o
    .mData_mData_5_valid   (featureWidthConvert_1_mData_mData_5_valid         ), //o
    .mData_mData_5_payload (featureWidthConvert_1_mData_mData_5_payload[127:0]), //o
    .mData_mData_6_valid   (featureWidthConvert_1_mData_mData_6_valid         ), //o
    .mData_mData_6_payload (featureWidthConvert_1_mData_mData_6_payload[127:0]), //o
    .mData_mData_7_valid   (featureWidthConvert_1_mData_mData_7_valid         ), //o
    .mData_mData_7_payload (featureWidthConvert_1_mData_mData_7_payload[127:0]), //o
    .mData_mData_8_valid   (featureWidthConvert_1_mData_mData_8_valid         ), //o
    .mData_mData_8_payload (featureWidthConvert_1_mData_mData_8_payload[127:0]), //o
    .mData_ready           (featureWidthConvert_1_mData_ready                 ), //i
    .rowNumIn              (rowNumIn[9:0]                                     ), //i
    .colNumIn              (colNumIn[9:0]                                     ), //i
    .start                 (featureWidthConvert_1_start                       ), //i
    .channelIn             (channelIn[11:0]                                   ), //i
    .reset                 (reset                                             ), //i
    .clk                   (clk                                               ), //i
    .softReset             (softReset                                         )  //i
  );
  FeatureConv11Convert featureConv11Convert_1 (
    .io_sData_valid           (featureConv11Convert_1_io_sData_valid                 ), //i
    .io_sData_ready           (featureConv11Convert_1_io_sData_ready                 ), //o
    .io_sData_payload         (featureConv11Convert_1_io_sData_payload[127:0]        ), //i
    .io_mData_mData_0_valid   (featureConv11Convert_1_io_mData_mData_0_valid         ), //o
    .io_mData_mData_0_payload (featureConv11Convert_1_io_mData_mData_0_payload[127:0]), //o
    .io_mData_mData_1_valid   (featureConv11Convert_1_io_mData_mData_1_valid         ), //o
    .io_mData_mData_1_payload (featureConv11Convert_1_io_mData_mData_1_payload[127:0]), //o
    .io_mData_mData_2_valid   (featureConv11Convert_1_io_mData_mData_2_valid         ), //o
    .io_mData_mData_2_payload (featureConv11Convert_1_io_mData_mData_2_payload[127:0]), //o
    .io_mData_mData_3_valid   (featureConv11Convert_1_io_mData_mData_3_valid         ), //o
    .io_mData_mData_3_payload (featureConv11Convert_1_io_mData_mData_3_payload[127:0]), //o
    .io_mData_mData_4_valid   (featureConv11Convert_1_io_mData_mData_4_valid         ), //o
    .io_mData_mData_4_payload (featureConv11Convert_1_io_mData_mData_4_payload[127:0]), //o
    .io_mData_mData_5_valid   (featureConv11Convert_1_io_mData_mData_5_valid         ), //o
    .io_mData_mData_5_payload (featureConv11Convert_1_io_mData_mData_5_payload[127:0]), //o
    .io_mData_mData_6_valid   (featureConv11Convert_1_io_mData_mData_6_valid         ), //o
    .io_mData_mData_6_payload (featureConv11Convert_1_io_mData_mData_6_payload[127:0]), //o
    .io_mData_mData_7_valid   (featureConv11Convert_1_io_mData_mData_7_valid         ), //o
    .io_mData_mData_7_payload (featureConv11Convert_1_io_mData_mData_7_payload[127:0]), //o
    .io_mData_mData_8_valid   (featureConv11Convert_1_io_mData_mData_8_valid         ), //o
    .io_mData_mData_8_payload (featureConv11Convert_1_io_mData_mData_8_payload[127:0]), //o
    .io_mData_ready           (featureConv11Convert_1_io_mData_ready                 ), //i
    .io_rowNumIn              (rowNumIn[9:0]                                         ), //i
    .io_colNumIn              (colNumIn[9:0]                                         ), //i
    .io_start                 (featureConv11Convert_1_io_start                       ), //i
    .io_channelIn             (channelIn[11:0]                                       ), //i
    .clk                      (clk                                                   ), //i
    .reset                    (reset                                                 ), //i
    .softReset                (softReset                                             )  //i
  );
  always @(*) begin
    case(convType)
      2'b00 : begin
        padding_1_sData_valid = sData_valid;
      end
      2'b01 : begin
        padding_1_sData_valid = 1'b0;
      end
      2'b10 : begin
        padding_1_sData_valid = 1'b0;
      end
      default : begin
        padding_1_sData_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        sData_ready = padding_1_sData_ready;
      end
      2'b01 : begin
        sData_ready = featureWidthConvert_1_sData_ready;
      end
      2'b10 : begin
        sData_ready = featureConv11Convert_1_io_sData_ready;
      end
      default : begin
        sData_ready = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        padding_1_sData_payload = sData_payload;
      end
      2'b01 : begin
        padding_1_sData_payload = 128'h0;
      end
      2'b10 : begin
        padding_1_sData_payload = 128'h0;
      end
      default : begin
        padding_1_sData_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        padding_1_start = start;
      end
      2'b01 : begin
        padding_1_start = 1'b0;
      end
      2'b10 : begin
        padding_1_start = 1'b0;
      end
      default : begin
        padding_1_start = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_0_valid = featureGenerate_1_mData_mData_0_valid;
      end
      2'b01 : begin
        mData_mData_0_valid = featureWidthConvert_1_mData_mData_0_valid;
      end
      2'b10 : begin
        mData_mData_0_valid = featureConv11Convert_1_io_mData_mData_0_valid;
      end
      default : begin
        mData_mData_0_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_0_payload = featureGenerate_1_mData_mData_0_payload;
      end
      2'b01 : begin
        mData_mData_0_payload = featureWidthConvert_1_mData_mData_0_payload;
      end
      2'b10 : begin
        mData_mData_0_payload = featureConv11Convert_1_io_mData_mData_0_payload;
      end
      default : begin
        mData_mData_0_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_1_valid = featureGenerate_1_mData_mData_1_valid;
      end
      2'b01 : begin
        mData_mData_1_valid = featureWidthConvert_1_mData_mData_1_valid;
      end
      2'b10 : begin
        mData_mData_1_valid = featureConv11Convert_1_io_mData_mData_1_valid;
      end
      default : begin
        mData_mData_1_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_1_payload = featureGenerate_1_mData_mData_1_payload;
      end
      2'b01 : begin
        mData_mData_1_payload = featureWidthConvert_1_mData_mData_1_payload;
      end
      2'b10 : begin
        mData_mData_1_payload = featureConv11Convert_1_io_mData_mData_1_payload;
      end
      default : begin
        mData_mData_1_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_2_valid = featureGenerate_1_mData_mData_2_valid;
      end
      2'b01 : begin
        mData_mData_2_valid = featureWidthConvert_1_mData_mData_2_valid;
      end
      2'b10 : begin
        mData_mData_2_valid = featureConv11Convert_1_io_mData_mData_2_valid;
      end
      default : begin
        mData_mData_2_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_2_payload = featureGenerate_1_mData_mData_2_payload;
      end
      2'b01 : begin
        mData_mData_2_payload = featureWidthConvert_1_mData_mData_2_payload;
      end
      2'b10 : begin
        mData_mData_2_payload = featureConv11Convert_1_io_mData_mData_2_payload;
      end
      default : begin
        mData_mData_2_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_3_valid = featureGenerate_1_mData_mData_3_valid;
      end
      2'b01 : begin
        mData_mData_3_valid = featureWidthConvert_1_mData_mData_3_valid;
      end
      2'b10 : begin
        mData_mData_3_valid = featureConv11Convert_1_io_mData_mData_3_valid;
      end
      default : begin
        mData_mData_3_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_3_payload = featureGenerate_1_mData_mData_3_payload;
      end
      2'b01 : begin
        mData_mData_3_payload = featureWidthConvert_1_mData_mData_3_payload;
      end
      2'b10 : begin
        mData_mData_3_payload = featureConv11Convert_1_io_mData_mData_3_payload;
      end
      default : begin
        mData_mData_3_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_4_valid = featureGenerate_1_mData_mData_4_valid;
      end
      2'b01 : begin
        mData_mData_4_valid = featureWidthConvert_1_mData_mData_4_valid;
      end
      2'b10 : begin
        mData_mData_4_valid = featureConv11Convert_1_io_mData_mData_4_valid;
      end
      default : begin
        mData_mData_4_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_4_payload = featureGenerate_1_mData_mData_4_payload;
      end
      2'b01 : begin
        mData_mData_4_payload = featureWidthConvert_1_mData_mData_4_payload;
      end
      2'b10 : begin
        mData_mData_4_payload = featureConv11Convert_1_io_mData_mData_4_payload;
      end
      default : begin
        mData_mData_4_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_5_valid = featureGenerate_1_mData_mData_5_valid;
      end
      2'b01 : begin
        mData_mData_5_valid = featureWidthConvert_1_mData_mData_5_valid;
      end
      2'b10 : begin
        mData_mData_5_valid = featureConv11Convert_1_io_mData_mData_5_valid;
      end
      default : begin
        mData_mData_5_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_5_payload = featureGenerate_1_mData_mData_5_payload;
      end
      2'b01 : begin
        mData_mData_5_payload = featureWidthConvert_1_mData_mData_5_payload;
      end
      2'b10 : begin
        mData_mData_5_payload = featureConv11Convert_1_io_mData_mData_5_payload;
      end
      default : begin
        mData_mData_5_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_6_valid = featureGenerate_1_mData_mData_6_valid;
      end
      2'b01 : begin
        mData_mData_6_valid = featureWidthConvert_1_mData_mData_6_valid;
      end
      2'b10 : begin
        mData_mData_6_valid = featureConv11Convert_1_io_mData_mData_6_valid;
      end
      default : begin
        mData_mData_6_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_6_payload = featureGenerate_1_mData_mData_6_payload;
      end
      2'b01 : begin
        mData_mData_6_payload = featureWidthConvert_1_mData_mData_6_payload;
      end
      2'b10 : begin
        mData_mData_6_payload = featureConv11Convert_1_io_mData_mData_6_payload;
      end
      default : begin
        mData_mData_6_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_7_valid = featureGenerate_1_mData_mData_7_valid;
      end
      2'b01 : begin
        mData_mData_7_valid = featureWidthConvert_1_mData_mData_7_valid;
      end
      2'b10 : begin
        mData_mData_7_valid = featureConv11Convert_1_io_mData_mData_7_valid;
      end
      default : begin
        mData_mData_7_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_7_payload = featureGenerate_1_mData_mData_7_payload;
      end
      2'b01 : begin
        mData_mData_7_payload = featureWidthConvert_1_mData_mData_7_payload;
      end
      2'b10 : begin
        mData_mData_7_payload = featureConv11Convert_1_io_mData_mData_7_payload;
      end
      default : begin
        mData_mData_7_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_8_valid = featureGenerate_1_mData_mData_8_valid;
      end
      2'b01 : begin
        mData_mData_8_valid = featureWidthConvert_1_mData_mData_8_valid;
      end
      2'b10 : begin
        mData_mData_8_valid = featureConv11Convert_1_io_mData_mData_8_valid;
      end
      default : begin
        mData_mData_8_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        mData_mData_8_payload = featureGenerate_1_mData_mData_8_payload;
      end
      2'b01 : begin
        mData_mData_8_payload = featureWidthConvert_1_mData_mData_8_payload;
      end
      2'b10 : begin
        mData_mData_8_payload = featureConv11Convert_1_io_mData_mData_8_payload;
      end
      default : begin
        mData_mData_8_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureGenerate_1_mData_ready = mData_ready;
      end
      2'b01 : begin
        featureGenerate_1_mData_ready = 1'b0;
      end
      2'b10 : begin
        featureGenerate_1_mData_ready = 1'b0;
      end
      default : begin
        featureGenerate_1_mData_ready = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureWidthConvert_1_sData_valid = 1'b0;
      end
      2'b01 : begin
        featureWidthConvert_1_sData_valid = sData_valid;
      end
      2'b10 : begin
        featureWidthConvert_1_sData_valid = 1'b0;
      end
      default : begin
        featureWidthConvert_1_sData_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureWidthConvert_1_sData_payload = 128'h0;
      end
      2'b01 : begin
        featureWidthConvert_1_sData_payload = sData_payload;
      end
      2'b10 : begin
        featureWidthConvert_1_sData_payload = 128'h0;
      end
      default : begin
        featureWidthConvert_1_sData_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureWidthConvert_1_mData_ready = 1'b0;
      end
      2'b01 : begin
        featureWidthConvert_1_mData_ready = mData_ready;
      end
      2'b10 : begin
        featureWidthConvert_1_mData_ready = 1'b0;
      end
      default : begin
        featureWidthConvert_1_mData_ready = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureWidthConvert_1_start = 1'b0;
      end
      2'b01 : begin
        featureWidthConvert_1_start = start;
      end
      2'b10 : begin
        featureWidthConvert_1_start = 1'b0;
      end
      default : begin
        featureWidthConvert_1_start = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureConv11Convert_1_io_sData_valid = 1'b0;
      end
      2'b01 : begin
        featureConv11Convert_1_io_sData_valid = 1'b0;
      end
      2'b10 : begin
        featureConv11Convert_1_io_sData_valid = sData_valid;
      end
      default : begin
        featureConv11Convert_1_io_sData_valid = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureConv11Convert_1_io_sData_payload = 128'h0;
      end
      2'b01 : begin
        featureConv11Convert_1_io_sData_payload = 128'h0;
      end
      2'b10 : begin
        featureConv11Convert_1_io_sData_payload = sData_payload;
      end
      default : begin
        featureConv11Convert_1_io_sData_payload = 128'h0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureConv11Convert_1_io_mData_ready = 1'b0;
      end
      2'b01 : begin
        featureConv11Convert_1_io_mData_ready = 1'b0;
      end
      2'b10 : begin
        featureConv11Convert_1_io_mData_ready = mData_ready;
      end
      default : begin
        featureConv11Convert_1_io_mData_ready = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(convType)
      2'b00 : begin
        featureConv11Convert_1_io_start = 1'b0;
      end
      2'b01 : begin
        featureConv11Convert_1_io_start = 1'b0;
      end
      2'b10 : begin
        featureConv11Convert_1_io_start = start;
      end
      default : begin
        featureConv11Convert_1_io_start = 1'b0;
      end
    endcase
  end


endmodule

module ChannelIncr (
  input               sData_valid,
  output              sData_ready,
  input      [7:0]    sData_payload,
  output              mData_valid,
  input               mData_ready,
  output     [127:0]  mData_payload
);


  assign sData_ready = mData_ready;
  assign mData_valid = sData_valid;
  assign mData_payload = {120'd0, sData_payload};

endmodule

module WaStreamFifoPipe (
  input               push_valid,
  output              push_ready,
  input      [127:0]  push_payload,
  output              pop_valid,
  input               pop_ready,
  output     [127:0]  pop_payload,
  input               flush,
  output     [14:0]   availability,
  input               clk,
  input               reset,
  input               softReset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [127:0]  fifo_io_pop_payload;
  wire       [14:0]   fifo_io_availability;
  reg        [127:0]  dataReg;
  wire                fifo_io_pop_fire;
  reg                 fireReg;
  reg                 validHold;
  wire                when_WaStreamFifoPipe_l26;
  reg        [127:0]  dataHold;
  wire                when_WaStreamFifoPipe_l30;

  StreamFifo fifo (
    .io_push_valid   (push_valid                ), //i
    .io_push_ready   (fifo_io_push_ready        ), //o
    .io_push_payload (push_payload[127:0]       ), //i
    .io_pop_valid    (fifo_io_pop_valid         ), //o
    .io_pop_ready    (pop_ready                 ), //i
    .io_pop_payload  (fifo_io_pop_payload[127:0]), //o
    .io_flush        (flush                     ), //i
    .io_availability (fifo_io_availability[14:0]), //o
    .clk             (clk                       ), //i
    .reset           (reset                     ), //i
    .softReset       (softReset                 )  //i
  );
  assign push_ready = fifo_io_push_ready;
  assign availability = fifo_io_availability;
  assign fifo_io_pop_fire = (fifo_io_pop_valid && pop_ready);
  assign when_WaStreamFifoPipe_l26 = (fireReg && (! pop_ready));
  assign when_WaStreamFifoPipe_l30 = (fireReg && (! pop_ready));
  assign pop_valid = (validHold || fireReg);
  assign pop_payload = (validHold ? dataHold : dataReg);
  always @(posedge clk) begin
    dataReg <= fifo_io_pop_payload;
    if(when_WaStreamFifoPipe_l26) begin
      dataHold <= dataReg;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      fireReg <= 1'b0;
      validHold <= 1'b0;
    end else begin
      if(softReset) begin
      fireReg <= 1'b0;
      validHold <= 1'b0;
      end else begin
        fireReg <= fifo_io_pop_fire;
        if(pop_ready) begin
          validHold <= 1'b0;
        end else begin
          if(when_WaStreamFifoPipe_l30) begin
            validHold <= 1'b1;
          end
        end
      end
    end
  end


endmodule

module LeakyRelu (
  input      [7:0]    dataIn_0,
  input      [7:0]    dataIn_1,
  input      [7:0]    dataIn_2,
  input      [7:0]    dataIn_3,
  input      [7:0]    dataIn_4,
  input      [7:0]    dataIn_5,
  input      [7:0]    dataIn_6,
  input      [7:0]    dataIn_7,
  input      [7:0]    dataIn_8,
  input      [7:0]    dataIn_9,
  input      [7:0]    dataIn_10,
  input      [7:0]    dataIn_11,
  input      [7:0]    dataIn_12,
  input      [7:0]    dataIn_13,
  input      [7:0]    dataIn_14,
  input      [7:0]    dataIn_15,
  input      [7:0]    quanZero,
  input      [31:0]   amendReg,
  output     [7:0]    dataOut_0,
  output     [7:0]    dataOut_1,
  output     [7:0]    dataOut_2,
  output     [7:0]    dataOut_3,
  output     [7:0]    dataOut_4,
  output     [7:0]    dataOut_5,
  output     [7:0]    dataOut_6,
  output     [7:0]    dataOut_7,
  output     [7:0]    dataOut_8,
  output     [7:0]    dataOut_9,
  output     [7:0]    dataOut_10,
  output     [7:0]    dataOut_11,
  output     [7:0]    dataOut_12,
  output     [7:0]    dataOut_13,
  output     [7:0]    dataOut_14,
  output     [7:0]    dataOut_15,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [15:0]   addSub_A;
  wire       [15:0]   addSub_2_A;
  wire       [15:0]   addSub_4_A;
  wire       [15:0]   addSub_6_A;
  wire       [15:0]   addSub_8_A;
  wire       [15:0]   addSub_10_A;
  wire       [15:0]   addSub_12_A;
  wire       [15:0]   addSub_14_A;
  wire       [15:0]   addSub_16_A;
  wire       [15:0]   addSub_18_A;
  wire       [15:0]   addSub_20_A;
  wire       [15:0]   addSub_22_A;
  wire       [15:0]   addSub_24_A;
  wire       [15:0]   addSub_26_A;
  wire       [15:0]   addSub_28_A;
  wire       [15:0]   addSub_30_A;
  wire       [15:0]   addSub_S;
  wire       [31:0]   mul_P;
  wire       [15:0]   addSub_1_S;
  wire       [15:0]   addSub_2_S;
  wire       [31:0]   mul_1_P;
  wire       [15:0]   addSub_3_S;
  wire       [15:0]   addSub_4_S;
  wire       [31:0]   mul_2_P;
  wire       [15:0]   addSub_5_S;
  wire       [15:0]   addSub_6_S;
  wire       [31:0]   mul_3_P;
  wire       [15:0]   addSub_7_S;
  wire       [15:0]   addSub_8_S;
  wire       [31:0]   mul_4_P;
  wire       [15:0]   addSub_9_S;
  wire       [15:0]   addSub_10_S;
  wire       [31:0]   mul_5_P;
  wire       [15:0]   addSub_11_S;
  wire       [15:0]   addSub_12_S;
  wire       [31:0]   mul_6_P;
  wire       [15:0]   addSub_13_S;
  wire       [15:0]   addSub_14_S;
  wire       [31:0]   mul_7_P;
  wire       [15:0]   addSub_15_S;
  wire       [15:0]   addSub_16_S;
  wire       [31:0]   mul_8_P;
  wire       [15:0]   addSub_17_S;
  wire       [15:0]   addSub_18_S;
  wire       [31:0]   mul_9_P;
  wire       [15:0]   addSub_19_S;
  wire       [15:0]   addSub_20_S;
  wire       [31:0]   mul_10_P;
  wire       [15:0]   addSub_21_S;
  wire       [15:0]   addSub_22_S;
  wire       [31:0]   mul_11_P;
  wire       [15:0]   addSub_23_S;
  wire       [15:0]   addSub_24_S;
  wire       [31:0]   mul_12_P;
  wire       [15:0]   addSub_25_S;
  wire       [15:0]   addSub_26_S;
  wire       [31:0]   mul_13_P;
  wire       [15:0]   addSub_27_S;
  wire       [15:0]   addSub_28_S;
  wire       [31:0]   mul_14_P;
  wire       [15:0]   addSub_29_S;
  wire       [15:0]   addSub_30_S;
  wire       [31:0]   mul_15_P;
  wire       [15:0]   addSub_31_S;
  wire       [14:0]   _zz__zz_A_1;
  wire       [14:0]   _zz__zz_A_1_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_32;
  wire       [15:0]   _zz_1;
  wire       [15:0]   _zz_2;
  wire       [15:0]   _zz_3;
  wire       [15:0]   _zz_4;
  wire       [15:0]   _zz_5;
  wire       [15:0]   _zz_6;
  wire       [15:0]   _zz_7;
  wire       [15:0]   _zz_8;
  wire       [15:0]   _zz_9;
  wire       [15:0]   _zz_10;
  wire       [15:0]   _zz_11;
  wire       [15:0]   _zz_12;
  wire       [15:0]   _zz_13;
  wire       [15:0]   _zz_14;
  wire       [15:0]   _zz_15;
  wire       [15:0]   _zz_16;
  wire       [15:0]   _zz__zz_A_3;
  wire       [15:0]   _zz__zz_A_3_1;
  wire       [15:0]   _zz__zz_A_3_2;
  wire       [15:0]   _zz__zz_A_3_3;
  wire       [15:0]   _zz__zz_A_3_4;
  wire       [15:0]   _zz__zz_A_3_5;
  wire       [15:0]   _zz__zz_A_3_6;
  wire       [15:0]   _zz__zz_A_3_7;
  wire       [15:0]   _zz__zz_A_3_8;
  wire       [15:0]   _zz__zz_A_3_9;
  wire       [15:0]   _zz__zz_A_3_10;
  wire       [15:0]   _zz__zz_A_3_11;
  wire       [15:0]   _zz__zz_A_3_12;
  wire       [15:0]   _zz__zz_A_3_13;
  wire       [15:0]   _zz__zz_A_3_14;
  wire       [15:0]   _zz__zz_A_3_15;
  wire       [15:0]   _zz__zz_A_3_16;
  wire       [15:0]   _zz__zz_A_3_17;
  wire       [15:0]   _zz__zz_A_3_18;
  wire       [15:0]   _zz__zz_A_3_19;
  wire       [15:0]   _zz__zz_A_3_20;
  wire       [15:0]   _zz__zz_A_3_21;
  wire       [15:0]   _zz__zz_A_3_22;
  wire       [15:0]   _zz__zz_A_3_23;
  wire       [15:0]   _zz__zz_A_3_24;
  wire       [15:0]   _zz__zz_A_3_25;
  wire       [15:0]   _zz__zz_A_3_26;
  wire       [15:0]   _zz__zz_A_3_27;
  wire       [15:0]   _zz__zz_A_3_28;
  wire       [15:0]   _zz__zz_A_3_29;
  wire       [15:0]   _zz__zz_A_3_30;
  wire       [15:0]   _zz__zz_A_3_31;
  wire       [15:0]   _zz__zz_dataOut_0;
  wire       [15:0]   _zz_when_LeakyRelu_l157;
  wire       [14:0]   _zz__zz_A_5;
  wire       [14:0]   _zz__zz_A_5_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_1_1;
  wire       [15:0]   _zz_17;
  wire       [15:0]   _zz_18;
  wire       [15:0]   _zz_19;
  wire       [15:0]   _zz_20;
  wire       [15:0]   _zz_21;
  wire       [15:0]   _zz_22;
  wire       [15:0]   _zz_23;
  wire       [15:0]   _zz_24;
  wire       [15:0]   _zz_25;
  wire       [15:0]   _zz_26;
  wire       [15:0]   _zz_27;
  wire       [15:0]   _zz_28;
  wire       [15:0]   _zz_29;
  wire       [15:0]   _zz_30;
  wire       [15:0]   _zz_31;
  wire       [15:0]   _zz_32;
  wire       [15:0]   _zz__zz_A_7;
  wire       [15:0]   _zz__zz_A_7_1;
  wire       [15:0]   _zz__zz_A_7_2;
  wire       [15:0]   _zz__zz_A_7_3;
  wire       [15:0]   _zz__zz_A_7_4;
  wire       [15:0]   _zz__zz_A_7_5;
  wire       [15:0]   _zz__zz_A_7_6;
  wire       [15:0]   _zz__zz_A_7_7;
  wire       [15:0]   _zz__zz_A_7_8;
  wire       [15:0]   _zz__zz_A_7_9;
  wire       [15:0]   _zz__zz_A_7_10;
  wire       [15:0]   _zz__zz_A_7_11;
  wire       [15:0]   _zz__zz_A_7_12;
  wire       [15:0]   _zz__zz_A_7_13;
  wire       [15:0]   _zz__zz_A_7_14;
  wire       [15:0]   _zz__zz_A_7_15;
  wire       [15:0]   _zz__zz_A_7_16;
  wire       [15:0]   _zz__zz_A_7_17;
  wire       [15:0]   _zz__zz_A_7_18;
  wire       [15:0]   _zz__zz_A_7_19;
  wire       [15:0]   _zz__zz_A_7_20;
  wire       [15:0]   _zz__zz_A_7_21;
  wire       [15:0]   _zz__zz_A_7_22;
  wire       [15:0]   _zz__zz_A_7_23;
  wire       [15:0]   _zz__zz_A_7_24;
  wire       [15:0]   _zz__zz_A_7_25;
  wire       [15:0]   _zz__zz_A_7_26;
  wire       [15:0]   _zz__zz_A_7_27;
  wire       [15:0]   _zz__zz_A_7_28;
  wire       [15:0]   _zz__zz_A_7_29;
  wire       [15:0]   _zz__zz_A_7_30;
  wire       [15:0]   _zz__zz_A_7_31;
  wire       [15:0]   _zz__zz_dataOut_1;
  wire       [15:0]   _zz_when_LeakyRelu_l157_1;
  wire       [14:0]   _zz__zz_A_9;
  wire       [14:0]   _zz__zz_A_9_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_2_1;
  wire       [15:0]   _zz_33;
  wire       [15:0]   _zz_34;
  wire       [15:0]   _zz_35;
  wire       [15:0]   _zz_36;
  wire       [15:0]   _zz_37;
  wire       [15:0]   _zz_38;
  wire       [15:0]   _zz_39;
  wire       [15:0]   _zz_40;
  wire       [15:0]   _zz_41;
  wire       [15:0]   _zz_42;
  wire       [15:0]   _zz_43;
  wire       [15:0]   _zz_44;
  wire       [15:0]   _zz_45;
  wire       [15:0]   _zz_46;
  wire       [15:0]   _zz_47;
  wire       [15:0]   _zz_48;
  wire       [15:0]   _zz__zz_A_11;
  wire       [15:0]   _zz__zz_A_11_1;
  wire       [15:0]   _zz__zz_A_11_2;
  wire       [15:0]   _zz__zz_A_11_3;
  wire       [15:0]   _zz__zz_A_11_4;
  wire       [15:0]   _zz__zz_A_11_5;
  wire       [15:0]   _zz__zz_A_11_6;
  wire       [15:0]   _zz__zz_A_11_7;
  wire       [15:0]   _zz__zz_A_11_8;
  wire       [15:0]   _zz__zz_A_11_9;
  wire       [15:0]   _zz__zz_A_11_10;
  wire       [15:0]   _zz__zz_A_11_11;
  wire       [15:0]   _zz__zz_A_11_12;
  wire       [15:0]   _zz__zz_A_11_13;
  wire       [15:0]   _zz__zz_A_11_14;
  wire       [15:0]   _zz__zz_A_11_15;
  wire       [15:0]   _zz__zz_A_11_16;
  wire       [15:0]   _zz__zz_A_11_17;
  wire       [15:0]   _zz__zz_A_11_18;
  wire       [15:0]   _zz__zz_A_11_19;
  wire       [15:0]   _zz__zz_A_11_20;
  wire       [15:0]   _zz__zz_A_11_21;
  wire       [15:0]   _zz__zz_A_11_22;
  wire       [15:0]   _zz__zz_A_11_23;
  wire       [15:0]   _zz__zz_A_11_24;
  wire       [15:0]   _zz__zz_A_11_25;
  wire       [15:0]   _zz__zz_A_11_26;
  wire       [15:0]   _zz__zz_A_11_27;
  wire       [15:0]   _zz__zz_A_11_28;
  wire       [15:0]   _zz__zz_A_11_29;
  wire       [15:0]   _zz__zz_A_11_30;
  wire       [15:0]   _zz__zz_A_11_31;
  wire       [15:0]   _zz__zz_dataOut_2;
  wire       [15:0]   _zz_when_LeakyRelu_l157_2;
  wire       [14:0]   _zz__zz_A_13;
  wire       [14:0]   _zz__zz_A_13_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_3_1;
  wire       [15:0]   _zz_49;
  wire       [15:0]   _zz_50;
  wire       [15:0]   _zz_51;
  wire       [15:0]   _zz_52;
  wire       [15:0]   _zz_53;
  wire       [15:0]   _zz_54;
  wire       [15:0]   _zz_55;
  wire       [15:0]   _zz_56;
  wire       [15:0]   _zz_57;
  wire       [15:0]   _zz_58;
  wire       [15:0]   _zz_59;
  wire       [15:0]   _zz_60;
  wire       [15:0]   _zz_61;
  wire       [15:0]   _zz_62;
  wire       [15:0]   _zz_63;
  wire       [15:0]   _zz_64;
  wire       [15:0]   _zz__zz_A_15;
  wire       [15:0]   _zz__zz_A_15_1;
  wire       [15:0]   _zz__zz_A_15_2;
  wire       [15:0]   _zz__zz_A_15_3;
  wire       [15:0]   _zz__zz_A_15_4;
  wire       [15:0]   _zz__zz_A_15_5;
  wire       [15:0]   _zz__zz_A_15_6;
  wire       [15:0]   _zz__zz_A_15_7;
  wire       [15:0]   _zz__zz_A_15_8;
  wire       [15:0]   _zz__zz_A_15_9;
  wire       [15:0]   _zz__zz_A_15_10;
  wire       [15:0]   _zz__zz_A_15_11;
  wire       [15:0]   _zz__zz_A_15_12;
  wire       [15:0]   _zz__zz_A_15_13;
  wire       [15:0]   _zz__zz_A_15_14;
  wire       [15:0]   _zz__zz_A_15_15;
  wire       [15:0]   _zz__zz_A_15_16;
  wire       [15:0]   _zz__zz_A_15_17;
  wire       [15:0]   _zz__zz_A_15_18;
  wire       [15:0]   _zz__zz_A_15_19;
  wire       [15:0]   _zz__zz_A_15_20;
  wire       [15:0]   _zz__zz_A_15_21;
  wire       [15:0]   _zz__zz_A_15_22;
  wire       [15:0]   _zz__zz_A_15_23;
  wire       [15:0]   _zz__zz_A_15_24;
  wire       [15:0]   _zz__zz_A_15_25;
  wire       [15:0]   _zz__zz_A_15_26;
  wire       [15:0]   _zz__zz_A_15_27;
  wire       [15:0]   _zz__zz_A_15_28;
  wire       [15:0]   _zz__zz_A_15_29;
  wire       [15:0]   _zz__zz_A_15_30;
  wire       [15:0]   _zz__zz_A_15_31;
  wire       [15:0]   _zz__zz_dataOut_3;
  wire       [15:0]   _zz_when_LeakyRelu_l157_3;
  wire       [14:0]   _zz__zz_A_17;
  wire       [14:0]   _zz__zz_A_17_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_4_1;
  wire       [15:0]   _zz_65;
  wire       [15:0]   _zz_66;
  wire       [15:0]   _zz_67;
  wire       [15:0]   _zz_68;
  wire       [15:0]   _zz_69;
  wire       [15:0]   _zz_70;
  wire       [15:0]   _zz_71;
  wire       [15:0]   _zz_72;
  wire       [15:0]   _zz_73;
  wire       [15:0]   _zz_74;
  wire       [15:0]   _zz_75;
  wire       [15:0]   _zz_76;
  wire       [15:0]   _zz_77;
  wire       [15:0]   _zz_78;
  wire       [15:0]   _zz_79;
  wire       [15:0]   _zz_80;
  wire       [15:0]   _zz__zz_A_19;
  wire       [15:0]   _zz__zz_A_19_1;
  wire       [15:0]   _zz__zz_A_19_2;
  wire       [15:0]   _zz__zz_A_19_3;
  wire       [15:0]   _zz__zz_A_19_4;
  wire       [15:0]   _zz__zz_A_19_5;
  wire       [15:0]   _zz__zz_A_19_6;
  wire       [15:0]   _zz__zz_A_19_7;
  wire       [15:0]   _zz__zz_A_19_8;
  wire       [15:0]   _zz__zz_A_19_9;
  wire       [15:0]   _zz__zz_A_19_10;
  wire       [15:0]   _zz__zz_A_19_11;
  wire       [15:0]   _zz__zz_A_19_12;
  wire       [15:0]   _zz__zz_A_19_13;
  wire       [15:0]   _zz__zz_A_19_14;
  wire       [15:0]   _zz__zz_A_19_15;
  wire       [15:0]   _zz__zz_A_19_16;
  wire       [15:0]   _zz__zz_A_19_17;
  wire       [15:0]   _zz__zz_A_19_18;
  wire       [15:0]   _zz__zz_A_19_19;
  wire       [15:0]   _zz__zz_A_19_20;
  wire       [15:0]   _zz__zz_A_19_21;
  wire       [15:0]   _zz__zz_A_19_22;
  wire       [15:0]   _zz__zz_A_19_23;
  wire       [15:0]   _zz__zz_A_19_24;
  wire       [15:0]   _zz__zz_A_19_25;
  wire       [15:0]   _zz__zz_A_19_26;
  wire       [15:0]   _zz__zz_A_19_27;
  wire       [15:0]   _zz__zz_A_19_28;
  wire       [15:0]   _zz__zz_A_19_29;
  wire       [15:0]   _zz__zz_A_19_30;
  wire       [15:0]   _zz__zz_A_19_31;
  wire       [15:0]   _zz__zz_dataOut_4;
  wire       [15:0]   _zz_when_LeakyRelu_l157_4;
  wire       [14:0]   _zz__zz_A_21;
  wire       [14:0]   _zz__zz_A_21_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_5_1;
  wire       [15:0]   _zz_81;
  wire       [15:0]   _zz_82;
  wire       [15:0]   _zz_83;
  wire       [15:0]   _zz_84;
  wire       [15:0]   _zz_85;
  wire       [15:0]   _zz_86;
  wire       [15:0]   _zz_87;
  wire       [15:0]   _zz_88;
  wire       [15:0]   _zz_89;
  wire       [15:0]   _zz_90;
  wire       [15:0]   _zz_91;
  wire       [15:0]   _zz_92;
  wire       [15:0]   _zz_93;
  wire       [15:0]   _zz_94;
  wire       [15:0]   _zz_95;
  wire       [15:0]   _zz_96;
  wire       [15:0]   _zz__zz_A_23;
  wire       [15:0]   _zz__zz_A_23_1;
  wire       [15:0]   _zz__zz_A_23_2;
  wire       [15:0]   _zz__zz_A_23_3;
  wire       [15:0]   _zz__zz_A_23_4;
  wire       [15:0]   _zz__zz_A_23_5;
  wire       [15:0]   _zz__zz_A_23_6;
  wire       [15:0]   _zz__zz_A_23_7;
  wire       [15:0]   _zz__zz_A_23_8;
  wire       [15:0]   _zz__zz_A_23_9;
  wire       [15:0]   _zz__zz_A_23_10;
  wire       [15:0]   _zz__zz_A_23_11;
  wire       [15:0]   _zz__zz_A_23_12;
  wire       [15:0]   _zz__zz_A_23_13;
  wire       [15:0]   _zz__zz_A_23_14;
  wire       [15:0]   _zz__zz_A_23_15;
  wire       [15:0]   _zz__zz_A_23_16;
  wire       [15:0]   _zz__zz_A_23_17;
  wire       [15:0]   _zz__zz_A_23_18;
  wire       [15:0]   _zz__zz_A_23_19;
  wire       [15:0]   _zz__zz_A_23_20;
  wire       [15:0]   _zz__zz_A_23_21;
  wire       [15:0]   _zz__zz_A_23_22;
  wire       [15:0]   _zz__zz_A_23_23;
  wire       [15:0]   _zz__zz_A_23_24;
  wire       [15:0]   _zz__zz_A_23_25;
  wire       [15:0]   _zz__zz_A_23_26;
  wire       [15:0]   _zz__zz_A_23_27;
  wire       [15:0]   _zz__zz_A_23_28;
  wire       [15:0]   _zz__zz_A_23_29;
  wire       [15:0]   _zz__zz_A_23_30;
  wire       [15:0]   _zz__zz_A_23_31;
  wire       [15:0]   _zz__zz_dataOut_5;
  wire       [15:0]   _zz_when_LeakyRelu_l157_5;
  wire       [14:0]   _zz__zz_A_25;
  wire       [14:0]   _zz__zz_A_25_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_6_1;
  wire       [15:0]   _zz_97;
  wire       [15:0]   _zz_98;
  wire       [15:0]   _zz_99;
  wire       [15:0]   _zz_100;
  wire       [15:0]   _zz_101;
  wire       [15:0]   _zz_102;
  wire       [15:0]   _zz_103;
  wire       [15:0]   _zz_104;
  wire       [15:0]   _zz_105;
  wire       [15:0]   _zz_106;
  wire       [15:0]   _zz_107;
  wire       [15:0]   _zz_108;
  wire       [15:0]   _zz_109;
  wire       [15:0]   _zz_110;
  wire       [15:0]   _zz_111;
  wire       [15:0]   _zz_112;
  wire       [15:0]   _zz__zz_A_27;
  wire       [15:0]   _zz__zz_A_27_1;
  wire       [15:0]   _zz__zz_A_27_2;
  wire       [15:0]   _zz__zz_A_27_3;
  wire       [15:0]   _zz__zz_A_27_4;
  wire       [15:0]   _zz__zz_A_27_5;
  wire       [15:0]   _zz__zz_A_27_6;
  wire       [15:0]   _zz__zz_A_27_7;
  wire       [15:0]   _zz__zz_A_27_8;
  wire       [15:0]   _zz__zz_A_27_9;
  wire       [15:0]   _zz__zz_A_27_10;
  wire       [15:0]   _zz__zz_A_27_11;
  wire       [15:0]   _zz__zz_A_27_12;
  wire       [15:0]   _zz__zz_A_27_13;
  wire       [15:0]   _zz__zz_A_27_14;
  wire       [15:0]   _zz__zz_A_27_15;
  wire       [15:0]   _zz__zz_A_27_16;
  wire       [15:0]   _zz__zz_A_27_17;
  wire       [15:0]   _zz__zz_A_27_18;
  wire       [15:0]   _zz__zz_A_27_19;
  wire       [15:0]   _zz__zz_A_27_20;
  wire       [15:0]   _zz__zz_A_27_21;
  wire       [15:0]   _zz__zz_A_27_22;
  wire       [15:0]   _zz__zz_A_27_23;
  wire       [15:0]   _zz__zz_A_27_24;
  wire       [15:0]   _zz__zz_A_27_25;
  wire       [15:0]   _zz__zz_A_27_26;
  wire       [15:0]   _zz__zz_A_27_27;
  wire       [15:0]   _zz__zz_A_27_28;
  wire       [15:0]   _zz__zz_A_27_29;
  wire       [15:0]   _zz__zz_A_27_30;
  wire       [15:0]   _zz__zz_A_27_31;
  wire       [15:0]   _zz__zz_dataOut_6;
  wire       [15:0]   _zz_when_LeakyRelu_l157_6;
  wire       [14:0]   _zz__zz_A_29;
  wire       [14:0]   _zz__zz_A_29_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_7_1;
  wire       [15:0]   _zz_113;
  wire       [15:0]   _zz_114;
  wire       [15:0]   _zz_115;
  wire       [15:0]   _zz_116;
  wire       [15:0]   _zz_117;
  wire       [15:0]   _zz_118;
  wire       [15:0]   _zz_119;
  wire       [15:0]   _zz_120;
  wire       [15:0]   _zz_121;
  wire       [15:0]   _zz_122;
  wire       [15:0]   _zz_123;
  wire       [15:0]   _zz_124;
  wire       [15:0]   _zz_125;
  wire       [15:0]   _zz_126;
  wire       [15:0]   _zz_127;
  wire       [15:0]   _zz_128;
  wire       [15:0]   _zz__zz_A_31;
  wire       [15:0]   _zz__zz_A_31_1;
  wire       [15:0]   _zz__zz_A_31_2;
  wire       [15:0]   _zz__zz_A_31_3;
  wire       [15:0]   _zz__zz_A_31_4;
  wire       [15:0]   _zz__zz_A_31_5;
  wire       [15:0]   _zz__zz_A_31_6;
  wire       [15:0]   _zz__zz_A_31_7;
  wire       [15:0]   _zz__zz_A_31_8;
  wire       [15:0]   _zz__zz_A_31_9;
  wire       [15:0]   _zz__zz_A_31_10;
  wire       [15:0]   _zz__zz_A_31_11;
  wire       [15:0]   _zz__zz_A_31_12;
  wire       [15:0]   _zz__zz_A_31_13;
  wire       [15:0]   _zz__zz_A_31_14;
  wire       [15:0]   _zz__zz_A_31_15;
  wire       [15:0]   _zz__zz_A_31_16;
  wire       [15:0]   _zz__zz_A_31_17;
  wire       [15:0]   _zz__zz_A_31_18;
  wire       [15:0]   _zz__zz_A_31_19;
  wire       [15:0]   _zz__zz_A_31_20;
  wire       [15:0]   _zz__zz_A_31_21;
  wire       [15:0]   _zz__zz_A_31_22;
  wire       [15:0]   _zz__zz_A_31_23;
  wire       [15:0]   _zz__zz_A_31_24;
  wire       [15:0]   _zz__zz_A_31_25;
  wire       [15:0]   _zz__zz_A_31_26;
  wire       [15:0]   _zz__zz_A_31_27;
  wire       [15:0]   _zz__zz_A_31_28;
  wire       [15:0]   _zz__zz_A_31_29;
  wire       [15:0]   _zz__zz_A_31_30;
  wire       [15:0]   _zz__zz_A_31_31;
  wire       [15:0]   _zz__zz_dataOut_7;
  wire       [15:0]   _zz_when_LeakyRelu_l157_7;
  wire       [14:0]   _zz__zz_A_33;
  wire       [14:0]   _zz__zz_A_33_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_8_1;
  wire       [15:0]   _zz_129;
  wire       [15:0]   _zz_130;
  wire       [15:0]   _zz_131;
  wire       [15:0]   _zz_132;
  wire       [15:0]   _zz_133;
  wire       [15:0]   _zz_134;
  wire       [15:0]   _zz_135;
  wire       [15:0]   _zz_136;
  wire       [15:0]   _zz_137;
  wire       [15:0]   _zz_138;
  wire       [15:0]   _zz_139;
  wire       [15:0]   _zz_140;
  wire       [15:0]   _zz_141;
  wire       [15:0]   _zz_142;
  wire       [15:0]   _zz_143;
  wire       [15:0]   _zz_144;
  wire       [15:0]   _zz__zz_A_35;
  wire       [15:0]   _zz__zz_A_35_1;
  wire       [15:0]   _zz__zz_A_35_2;
  wire       [15:0]   _zz__zz_A_35_3;
  wire       [15:0]   _zz__zz_A_35_4;
  wire       [15:0]   _zz__zz_A_35_5;
  wire       [15:0]   _zz__zz_A_35_6;
  wire       [15:0]   _zz__zz_A_35_7;
  wire       [15:0]   _zz__zz_A_35_8;
  wire       [15:0]   _zz__zz_A_35_9;
  wire       [15:0]   _zz__zz_A_35_10;
  wire       [15:0]   _zz__zz_A_35_11;
  wire       [15:0]   _zz__zz_A_35_12;
  wire       [15:0]   _zz__zz_A_35_13;
  wire       [15:0]   _zz__zz_A_35_14;
  wire       [15:0]   _zz__zz_A_35_15;
  wire       [15:0]   _zz__zz_A_35_16;
  wire       [15:0]   _zz__zz_A_35_17;
  wire       [15:0]   _zz__zz_A_35_18;
  wire       [15:0]   _zz__zz_A_35_19;
  wire       [15:0]   _zz__zz_A_35_20;
  wire       [15:0]   _zz__zz_A_35_21;
  wire       [15:0]   _zz__zz_A_35_22;
  wire       [15:0]   _zz__zz_A_35_23;
  wire       [15:0]   _zz__zz_A_35_24;
  wire       [15:0]   _zz__zz_A_35_25;
  wire       [15:0]   _zz__zz_A_35_26;
  wire       [15:0]   _zz__zz_A_35_27;
  wire       [15:0]   _zz__zz_A_35_28;
  wire       [15:0]   _zz__zz_A_35_29;
  wire       [15:0]   _zz__zz_A_35_30;
  wire       [15:0]   _zz__zz_A_35_31;
  wire       [15:0]   _zz__zz_dataOut_8;
  wire       [15:0]   _zz_when_LeakyRelu_l157_8;
  wire       [14:0]   _zz__zz_A_37;
  wire       [14:0]   _zz__zz_A_37_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_9_1;
  wire       [15:0]   _zz_145;
  wire       [15:0]   _zz_146;
  wire       [15:0]   _zz_147;
  wire       [15:0]   _zz_148;
  wire       [15:0]   _zz_149;
  wire       [15:0]   _zz_150;
  wire       [15:0]   _zz_151;
  wire       [15:0]   _zz_152;
  wire       [15:0]   _zz_153;
  wire       [15:0]   _zz_154;
  wire       [15:0]   _zz_155;
  wire       [15:0]   _zz_156;
  wire       [15:0]   _zz_157;
  wire       [15:0]   _zz_158;
  wire       [15:0]   _zz_159;
  wire       [15:0]   _zz_160;
  wire       [15:0]   _zz__zz_A_39;
  wire       [15:0]   _zz__zz_A_39_1;
  wire       [15:0]   _zz__zz_A_39_2;
  wire       [15:0]   _zz__zz_A_39_3;
  wire       [15:0]   _zz__zz_A_39_4;
  wire       [15:0]   _zz__zz_A_39_5;
  wire       [15:0]   _zz__zz_A_39_6;
  wire       [15:0]   _zz__zz_A_39_7;
  wire       [15:0]   _zz__zz_A_39_8;
  wire       [15:0]   _zz__zz_A_39_9;
  wire       [15:0]   _zz__zz_A_39_10;
  wire       [15:0]   _zz__zz_A_39_11;
  wire       [15:0]   _zz__zz_A_39_12;
  wire       [15:0]   _zz__zz_A_39_13;
  wire       [15:0]   _zz__zz_A_39_14;
  wire       [15:0]   _zz__zz_A_39_15;
  wire       [15:0]   _zz__zz_A_39_16;
  wire       [15:0]   _zz__zz_A_39_17;
  wire       [15:0]   _zz__zz_A_39_18;
  wire       [15:0]   _zz__zz_A_39_19;
  wire       [15:0]   _zz__zz_A_39_20;
  wire       [15:0]   _zz__zz_A_39_21;
  wire       [15:0]   _zz__zz_A_39_22;
  wire       [15:0]   _zz__zz_A_39_23;
  wire       [15:0]   _zz__zz_A_39_24;
  wire       [15:0]   _zz__zz_A_39_25;
  wire       [15:0]   _zz__zz_A_39_26;
  wire       [15:0]   _zz__zz_A_39_27;
  wire       [15:0]   _zz__zz_A_39_28;
  wire       [15:0]   _zz__zz_A_39_29;
  wire       [15:0]   _zz__zz_A_39_30;
  wire       [15:0]   _zz__zz_A_39_31;
  wire       [15:0]   _zz__zz_dataOut_9;
  wire       [15:0]   _zz_when_LeakyRelu_l157_9;
  wire       [14:0]   _zz__zz_A_41;
  wire       [14:0]   _zz__zz_A_41_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_10_1;
  wire       [15:0]   _zz_161;
  wire       [15:0]   _zz_162;
  wire       [15:0]   _zz_163;
  wire       [15:0]   _zz_164;
  wire       [15:0]   _zz_165;
  wire       [15:0]   _zz_166;
  wire       [15:0]   _zz_167;
  wire       [15:0]   _zz_168;
  wire       [15:0]   _zz_169;
  wire       [15:0]   _zz_170;
  wire       [15:0]   _zz_171;
  wire       [15:0]   _zz_172;
  wire       [15:0]   _zz_173;
  wire       [15:0]   _zz_174;
  wire       [15:0]   _zz_175;
  wire       [15:0]   _zz_176;
  wire       [15:0]   _zz__zz_A_43;
  wire       [15:0]   _zz__zz_A_43_1;
  wire       [15:0]   _zz__zz_A_43_2;
  wire       [15:0]   _zz__zz_A_43_3;
  wire       [15:0]   _zz__zz_A_43_4;
  wire       [15:0]   _zz__zz_A_43_5;
  wire       [15:0]   _zz__zz_A_43_6;
  wire       [15:0]   _zz__zz_A_43_7;
  wire       [15:0]   _zz__zz_A_43_8;
  wire       [15:0]   _zz__zz_A_43_9;
  wire       [15:0]   _zz__zz_A_43_10;
  wire       [15:0]   _zz__zz_A_43_11;
  wire       [15:0]   _zz__zz_A_43_12;
  wire       [15:0]   _zz__zz_A_43_13;
  wire       [15:0]   _zz__zz_A_43_14;
  wire       [15:0]   _zz__zz_A_43_15;
  wire       [15:0]   _zz__zz_A_43_16;
  wire       [15:0]   _zz__zz_A_43_17;
  wire       [15:0]   _zz__zz_A_43_18;
  wire       [15:0]   _zz__zz_A_43_19;
  wire       [15:0]   _zz__zz_A_43_20;
  wire       [15:0]   _zz__zz_A_43_21;
  wire       [15:0]   _zz__zz_A_43_22;
  wire       [15:0]   _zz__zz_A_43_23;
  wire       [15:0]   _zz__zz_A_43_24;
  wire       [15:0]   _zz__zz_A_43_25;
  wire       [15:0]   _zz__zz_A_43_26;
  wire       [15:0]   _zz__zz_A_43_27;
  wire       [15:0]   _zz__zz_A_43_28;
  wire       [15:0]   _zz__zz_A_43_29;
  wire       [15:0]   _zz__zz_A_43_30;
  wire       [15:0]   _zz__zz_A_43_31;
  wire       [15:0]   _zz__zz_dataOut_10;
  wire       [15:0]   _zz_when_LeakyRelu_l157_10;
  wire       [14:0]   _zz__zz_A_45;
  wire       [14:0]   _zz__zz_A_45_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_11_1;
  wire       [15:0]   _zz_177;
  wire       [15:0]   _zz_178;
  wire       [15:0]   _zz_179;
  wire       [15:0]   _zz_180;
  wire       [15:0]   _zz_181;
  wire       [15:0]   _zz_182;
  wire       [15:0]   _zz_183;
  wire       [15:0]   _zz_184;
  wire       [15:0]   _zz_185;
  wire       [15:0]   _zz_186;
  wire       [15:0]   _zz_187;
  wire       [15:0]   _zz_188;
  wire       [15:0]   _zz_189;
  wire       [15:0]   _zz_190;
  wire       [15:0]   _zz_191;
  wire       [15:0]   _zz_192;
  wire       [15:0]   _zz__zz_A_47;
  wire       [15:0]   _zz__zz_A_47_1;
  wire       [15:0]   _zz__zz_A_47_2;
  wire       [15:0]   _zz__zz_A_47_3;
  wire       [15:0]   _zz__zz_A_47_4;
  wire       [15:0]   _zz__zz_A_47_5;
  wire       [15:0]   _zz__zz_A_47_6;
  wire       [15:0]   _zz__zz_A_47_7;
  wire       [15:0]   _zz__zz_A_47_8;
  wire       [15:0]   _zz__zz_A_47_9;
  wire       [15:0]   _zz__zz_A_47_10;
  wire       [15:0]   _zz__zz_A_47_11;
  wire       [15:0]   _zz__zz_A_47_12;
  wire       [15:0]   _zz__zz_A_47_13;
  wire       [15:0]   _zz__zz_A_47_14;
  wire       [15:0]   _zz__zz_A_47_15;
  wire       [15:0]   _zz__zz_A_47_16;
  wire       [15:0]   _zz__zz_A_47_17;
  wire       [15:0]   _zz__zz_A_47_18;
  wire       [15:0]   _zz__zz_A_47_19;
  wire       [15:0]   _zz__zz_A_47_20;
  wire       [15:0]   _zz__zz_A_47_21;
  wire       [15:0]   _zz__zz_A_47_22;
  wire       [15:0]   _zz__zz_A_47_23;
  wire       [15:0]   _zz__zz_A_47_24;
  wire       [15:0]   _zz__zz_A_47_25;
  wire       [15:0]   _zz__zz_A_47_26;
  wire       [15:0]   _zz__zz_A_47_27;
  wire       [15:0]   _zz__zz_A_47_28;
  wire       [15:0]   _zz__zz_A_47_29;
  wire       [15:0]   _zz__zz_A_47_30;
  wire       [15:0]   _zz__zz_A_47_31;
  wire       [15:0]   _zz__zz_dataOut_11;
  wire       [15:0]   _zz_when_LeakyRelu_l157_11;
  wire       [14:0]   _zz__zz_A_49;
  wire       [14:0]   _zz__zz_A_49_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_12_1;
  wire       [15:0]   _zz_193;
  wire       [15:0]   _zz_194;
  wire       [15:0]   _zz_195;
  wire       [15:0]   _zz_196;
  wire       [15:0]   _zz_197;
  wire       [15:0]   _zz_198;
  wire       [15:0]   _zz_199;
  wire       [15:0]   _zz_200;
  wire       [15:0]   _zz_201;
  wire       [15:0]   _zz_202;
  wire       [15:0]   _zz_203;
  wire       [15:0]   _zz_204;
  wire       [15:0]   _zz_205;
  wire       [15:0]   _zz_206;
  wire       [15:0]   _zz_207;
  wire       [15:0]   _zz_208;
  wire       [15:0]   _zz__zz_A_51;
  wire       [15:0]   _zz__zz_A_51_1;
  wire       [15:0]   _zz__zz_A_51_2;
  wire       [15:0]   _zz__zz_A_51_3;
  wire       [15:0]   _zz__zz_A_51_4;
  wire       [15:0]   _zz__zz_A_51_5;
  wire       [15:0]   _zz__zz_A_51_6;
  wire       [15:0]   _zz__zz_A_51_7;
  wire       [15:0]   _zz__zz_A_51_8;
  wire       [15:0]   _zz__zz_A_51_9;
  wire       [15:0]   _zz__zz_A_51_10;
  wire       [15:0]   _zz__zz_A_51_11;
  wire       [15:0]   _zz__zz_A_51_12;
  wire       [15:0]   _zz__zz_A_51_13;
  wire       [15:0]   _zz__zz_A_51_14;
  wire       [15:0]   _zz__zz_A_51_15;
  wire       [15:0]   _zz__zz_A_51_16;
  wire       [15:0]   _zz__zz_A_51_17;
  wire       [15:0]   _zz__zz_A_51_18;
  wire       [15:0]   _zz__zz_A_51_19;
  wire       [15:0]   _zz__zz_A_51_20;
  wire       [15:0]   _zz__zz_A_51_21;
  wire       [15:0]   _zz__zz_A_51_22;
  wire       [15:0]   _zz__zz_A_51_23;
  wire       [15:0]   _zz__zz_A_51_24;
  wire       [15:0]   _zz__zz_A_51_25;
  wire       [15:0]   _zz__zz_A_51_26;
  wire       [15:0]   _zz__zz_A_51_27;
  wire       [15:0]   _zz__zz_A_51_28;
  wire       [15:0]   _zz__zz_A_51_29;
  wire       [15:0]   _zz__zz_A_51_30;
  wire       [15:0]   _zz__zz_A_51_31;
  wire       [15:0]   _zz__zz_dataOut_12;
  wire       [15:0]   _zz_when_LeakyRelu_l157_12;
  wire       [14:0]   _zz__zz_A_53;
  wire       [14:0]   _zz__zz_A_53_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_13_1;
  wire       [15:0]   _zz_209;
  wire       [15:0]   _zz_210;
  wire       [15:0]   _zz_211;
  wire       [15:0]   _zz_212;
  wire       [15:0]   _zz_213;
  wire       [15:0]   _zz_214;
  wire       [15:0]   _zz_215;
  wire       [15:0]   _zz_216;
  wire       [15:0]   _zz_217;
  wire       [15:0]   _zz_218;
  wire       [15:0]   _zz_219;
  wire       [15:0]   _zz_220;
  wire       [15:0]   _zz_221;
  wire       [15:0]   _zz_222;
  wire       [15:0]   _zz_223;
  wire       [15:0]   _zz_224;
  wire       [15:0]   _zz__zz_A_55;
  wire       [15:0]   _zz__zz_A_55_1;
  wire       [15:0]   _zz__zz_A_55_2;
  wire       [15:0]   _zz__zz_A_55_3;
  wire       [15:0]   _zz__zz_A_55_4;
  wire       [15:0]   _zz__zz_A_55_5;
  wire       [15:0]   _zz__zz_A_55_6;
  wire       [15:0]   _zz__zz_A_55_7;
  wire       [15:0]   _zz__zz_A_55_8;
  wire       [15:0]   _zz__zz_A_55_9;
  wire       [15:0]   _zz__zz_A_55_10;
  wire       [15:0]   _zz__zz_A_55_11;
  wire       [15:0]   _zz__zz_A_55_12;
  wire       [15:0]   _zz__zz_A_55_13;
  wire       [15:0]   _zz__zz_A_55_14;
  wire       [15:0]   _zz__zz_A_55_15;
  wire       [15:0]   _zz__zz_A_55_16;
  wire       [15:0]   _zz__zz_A_55_17;
  wire       [15:0]   _zz__zz_A_55_18;
  wire       [15:0]   _zz__zz_A_55_19;
  wire       [15:0]   _zz__zz_A_55_20;
  wire       [15:0]   _zz__zz_A_55_21;
  wire       [15:0]   _zz__zz_A_55_22;
  wire       [15:0]   _zz__zz_A_55_23;
  wire       [15:0]   _zz__zz_A_55_24;
  wire       [15:0]   _zz__zz_A_55_25;
  wire       [15:0]   _zz__zz_A_55_26;
  wire       [15:0]   _zz__zz_A_55_27;
  wire       [15:0]   _zz__zz_A_55_28;
  wire       [15:0]   _zz__zz_A_55_29;
  wire       [15:0]   _zz__zz_A_55_30;
  wire       [15:0]   _zz__zz_A_55_31;
  wire       [15:0]   _zz__zz_dataOut_13;
  wire       [15:0]   _zz_when_LeakyRelu_l157_13;
  wire       [14:0]   _zz__zz_A_57;
  wire       [14:0]   _zz__zz_A_57_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_14_1;
  wire       [15:0]   _zz_225;
  wire       [15:0]   _zz_226;
  wire       [15:0]   _zz_227;
  wire       [15:0]   _zz_228;
  wire       [15:0]   _zz_229;
  wire       [15:0]   _zz_230;
  wire       [15:0]   _zz_231;
  wire       [15:0]   _zz_232;
  wire       [15:0]   _zz_233;
  wire       [15:0]   _zz_234;
  wire       [15:0]   _zz_235;
  wire       [15:0]   _zz_236;
  wire       [15:0]   _zz_237;
  wire       [15:0]   _zz_238;
  wire       [15:0]   _zz_239;
  wire       [15:0]   _zz_240;
  wire       [15:0]   _zz__zz_A_59;
  wire       [15:0]   _zz__zz_A_59_1;
  wire       [15:0]   _zz__zz_A_59_2;
  wire       [15:0]   _zz__zz_A_59_3;
  wire       [15:0]   _zz__zz_A_59_4;
  wire       [15:0]   _zz__zz_A_59_5;
  wire       [15:0]   _zz__zz_A_59_6;
  wire       [15:0]   _zz__zz_A_59_7;
  wire       [15:0]   _zz__zz_A_59_8;
  wire       [15:0]   _zz__zz_A_59_9;
  wire       [15:0]   _zz__zz_A_59_10;
  wire       [15:0]   _zz__zz_A_59_11;
  wire       [15:0]   _zz__zz_A_59_12;
  wire       [15:0]   _zz__zz_A_59_13;
  wire       [15:0]   _zz__zz_A_59_14;
  wire       [15:0]   _zz__zz_A_59_15;
  wire       [15:0]   _zz__zz_A_59_16;
  wire       [15:0]   _zz__zz_A_59_17;
  wire       [15:0]   _zz__zz_A_59_18;
  wire       [15:0]   _zz__zz_A_59_19;
  wire       [15:0]   _zz__zz_A_59_20;
  wire       [15:0]   _zz__zz_A_59_21;
  wire       [15:0]   _zz__zz_A_59_22;
  wire       [15:0]   _zz__zz_A_59_23;
  wire       [15:0]   _zz__zz_A_59_24;
  wire       [15:0]   _zz__zz_A_59_25;
  wire       [15:0]   _zz__zz_A_59_26;
  wire       [15:0]   _zz__zz_A_59_27;
  wire       [15:0]   _zz__zz_A_59_28;
  wire       [15:0]   _zz__zz_A_59_29;
  wire       [15:0]   _zz__zz_A_59_30;
  wire       [15:0]   _zz__zz_A_59_31;
  wire       [15:0]   _zz__zz_dataOut_14;
  wire       [15:0]   _zz_when_LeakyRelu_l157_14;
  wire       [14:0]   _zz__zz_A_61;
  wire       [14:0]   _zz__zz_A_61_1;
  wire       [3:0]    _zz_when_LeakyRelu_l101_15_1;
  wire       [15:0]   _zz_241;
  wire       [15:0]   _zz_242;
  wire       [15:0]   _zz_243;
  wire       [15:0]   _zz_244;
  wire       [15:0]   _zz_245;
  wire       [15:0]   _zz_246;
  wire       [15:0]   _zz_247;
  wire       [15:0]   _zz_248;
  wire       [15:0]   _zz_249;
  wire       [15:0]   _zz_250;
  wire       [15:0]   _zz_251;
  wire       [15:0]   _zz_252;
  wire       [15:0]   _zz_253;
  wire       [15:0]   _zz_254;
  wire       [15:0]   _zz_255;
  wire       [15:0]   _zz_256;
  wire       [15:0]   _zz__zz_A_63;
  wire       [15:0]   _zz__zz_A_63_1;
  wire       [15:0]   _zz__zz_A_63_2;
  wire       [15:0]   _zz__zz_A_63_3;
  wire       [15:0]   _zz__zz_A_63_4;
  wire       [15:0]   _zz__zz_A_63_5;
  wire       [15:0]   _zz__zz_A_63_6;
  wire       [15:0]   _zz__zz_A_63_7;
  wire       [15:0]   _zz__zz_A_63_8;
  wire       [15:0]   _zz__zz_A_63_9;
  wire       [15:0]   _zz__zz_A_63_10;
  wire       [15:0]   _zz__zz_A_63_11;
  wire       [15:0]   _zz__zz_A_63_12;
  wire       [15:0]   _zz__zz_A_63_13;
  wire       [15:0]   _zz__zz_A_63_14;
  wire       [15:0]   _zz__zz_A_63_15;
  wire       [15:0]   _zz__zz_A_63_16;
  wire       [15:0]   _zz__zz_A_63_17;
  wire       [15:0]   _zz__zz_A_63_18;
  wire       [15:0]   _zz__zz_A_63_19;
  wire       [15:0]   _zz__zz_A_63_20;
  wire       [15:0]   _zz__zz_A_63_21;
  wire       [15:0]   _zz__zz_A_63_22;
  wire       [15:0]   _zz__zz_A_63_23;
  wire       [15:0]   _zz__zz_A_63_24;
  wire       [15:0]   _zz__zz_A_63_25;
  wire       [15:0]   _zz__zz_A_63_26;
  wire       [15:0]   _zz__zz_A_63_27;
  wire       [15:0]   _zz__zz_A_63_28;
  wire       [15:0]   _zz__zz_A_63_29;
  wire       [15:0]   _zz__zz_A_63_30;
  wire       [15:0]   _zz__zz_A_63_31;
  wire       [15:0]   _zz__zz_dataOut_15;
  wire       [15:0]   _zz_when_LeakyRelu_l157_15;
  wire       [15:0]   leaky;
  reg        [7:0]    _zz_dataOut_0;
  reg        [15:0]   _zz_A;
  wire       [15:0]   _zz_when_LeakyRelu_l100;
  wire       [31:0]   _zz_when_LeakyRelu_l101;
  wire       [3:0]    _zz_when_LeakyRelu_l101_1;
  wire       [14:0]   _zz_A_1;
  wire       [14:0]   _zz_A_2;
  reg        [15:0]   _zz_when_LeakyRelu_l100_1;
  reg        [15:0]   _zz_when_LeakyRelu_l100_2;
  reg        [15:0]   _zz_when_LeakyRelu_l100_3;
  wire                when_LeakyRelu_l100;
  wire                when_LeakyRelu_l101;
  wire                when_LeakyRelu_l104;
  wire                when_LeakyRelu_l110;
  wire                when_LeakyRelu_l103;
  reg        [15:0]   _zz_A_3;
  reg        [15:0]   _zz_when_LeakyRelu_l100_3_regNext;
  wire                when_LeakyRelu_l127;
  wire                when_LeakyRelu_l131;
  wire                when_LeakyRelu_l133;
  wire                when_LeakyRelu_l131_1;
  wire                when_LeakyRelu_l133_1;
  wire                when_LeakyRelu_l131_2;
  wire                when_LeakyRelu_l133_2;
  wire                when_LeakyRelu_l131_3;
  wire                when_LeakyRelu_l133_3;
  wire                when_LeakyRelu_l131_4;
  wire                when_LeakyRelu_l133_4;
  wire                when_LeakyRelu_l131_5;
  wire                when_LeakyRelu_l133_5;
  wire                when_LeakyRelu_l131_6;
  wire                when_LeakyRelu_l133_6;
  wire                when_LeakyRelu_l131_7;
  wire                when_LeakyRelu_l133_7;
  wire                when_LeakyRelu_l131_8;
  wire                when_LeakyRelu_l133_8;
  wire                when_LeakyRelu_l131_9;
  wire                when_LeakyRelu_l133_9;
  wire                when_LeakyRelu_l131_10;
  wire                when_LeakyRelu_l133_10;
  wire                when_LeakyRelu_l131_11;
  wire                when_LeakyRelu_l133_11;
  wire                when_LeakyRelu_l131_12;
  wire                when_LeakyRelu_l133_12;
  wire                when_LeakyRelu_l131_13;
  wire                when_LeakyRelu_l133_13;
  wire                when_LeakyRelu_l131_14;
  wire                when_LeakyRelu_l133_14;
  wire                when_LeakyRelu_l131_15;
  wire                when_LeakyRelu_l133_15;
  wire       [15:0]   _zz_dataOut_0_1;
  wire                when_LeakyRelu_l155;
  wire                when_LeakyRelu_l157;
  reg        [7:0]    _zz_dataOut_1;
  reg        [15:0]   _zz_A_4;
  wire       [15:0]   _zz_when_LeakyRelu_l100_4;
  wire       [31:0]   _zz_when_LeakyRelu_l101_2;
  wire       [3:0]    _zz_when_LeakyRelu_l101_3;
  wire       [14:0]   _zz_A_5;
  wire       [14:0]   _zz_A_6;
  reg        [15:0]   _zz_when_LeakyRelu_l100_5;
  reg        [15:0]   _zz_when_LeakyRelu_l100_6;
  reg        [15:0]   _zz_when_LeakyRelu_l100_7;
  wire                when_LeakyRelu_l100_1;
  wire                when_LeakyRelu_l101_1;
  wire                when_LeakyRelu_l104_1;
  wire                when_LeakyRelu_l110_1;
  wire                when_LeakyRelu_l103_1;
  reg        [15:0]   _zz_A_7;
  reg        [15:0]   _zz_when_LeakyRelu_l100_7_regNext;
  wire                when_LeakyRelu_l127_1;
  wire                when_LeakyRelu_l131_16;
  wire                when_LeakyRelu_l133_16;
  wire                when_LeakyRelu_l131_17;
  wire                when_LeakyRelu_l133_17;
  wire                when_LeakyRelu_l131_18;
  wire                when_LeakyRelu_l133_18;
  wire                when_LeakyRelu_l131_19;
  wire                when_LeakyRelu_l133_19;
  wire                when_LeakyRelu_l131_20;
  wire                when_LeakyRelu_l133_20;
  wire                when_LeakyRelu_l131_21;
  wire                when_LeakyRelu_l133_21;
  wire                when_LeakyRelu_l131_22;
  wire                when_LeakyRelu_l133_22;
  wire                when_LeakyRelu_l131_23;
  wire                when_LeakyRelu_l133_23;
  wire                when_LeakyRelu_l131_24;
  wire                when_LeakyRelu_l133_24;
  wire                when_LeakyRelu_l131_25;
  wire                when_LeakyRelu_l133_25;
  wire                when_LeakyRelu_l131_26;
  wire                when_LeakyRelu_l133_26;
  wire                when_LeakyRelu_l131_27;
  wire                when_LeakyRelu_l133_27;
  wire                when_LeakyRelu_l131_28;
  wire                when_LeakyRelu_l133_28;
  wire                when_LeakyRelu_l131_29;
  wire                when_LeakyRelu_l133_29;
  wire                when_LeakyRelu_l131_30;
  wire                when_LeakyRelu_l133_30;
  wire                when_LeakyRelu_l131_31;
  wire                when_LeakyRelu_l133_31;
  wire       [15:0]   _zz_dataOut_1_1;
  wire                when_LeakyRelu_l155_1;
  wire                when_LeakyRelu_l157_1;
  reg        [7:0]    _zz_dataOut_2;
  reg        [15:0]   _zz_A_8;
  wire       [15:0]   _zz_when_LeakyRelu_l100_8;
  wire       [31:0]   _zz_when_LeakyRelu_l101_4;
  wire       [3:0]    _zz_when_LeakyRelu_l101_5;
  wire       [14:0]   _zz_A_9;
  wire       [14:0]   _zz_A_10;
  reg        [15:0]   _zz_when_LeakyRelu_l100_9;
  reg        [15:0]   _zz_when_LeakyRelu_l100_10;
  reg        [15:0]   _zz_when_LeakyRelu_l100_11;
  wire                when_LeakyRelu_l100_2;
  wire                when_LeakyRelu_l101_2;
  wire                when_LeakyRelu_l104_2;
  wire                when_LeakyRelu_l110_2;
  wire                when_LeakyRelu_l103_2;
  reg        [15:0]   _zz_A_11;
  reg        [15:0]   _zz_when_LeakyRelu_l100_11_regNext;
  wire                when_LeakyRelu_l127_2;
  wire                when_LeakyRelu_l131_32;
  wire                when_LeakyRelu_l133_32;
  wire                when_LeakyRelu_l131_33;
  wire                when_LeakyRelu_l133_33;
  wire                when_LeakyRelu_l131_34;
  wire                when_LeakyRelu_l133_34;
  wire                when_LeakyRelu_l131_35;
  wire                when_LeakyRelu_l133_35;
  wire                when_LeakyRelu_l131_36;
  wire                when_LeakyRelu_l133_36;
  wire                when_LeakyRelu_l131_37;
  wire                when_LeakyRelu_l133_37;
  wire                when_LeakyRelu_l131_38;
  wire                when_LeakyRelu_l133_38;
  wire                when_LeakyRelu_l131_39;
  wire                when_LeakyRelu_l133_39;
  wire                when_LeakyRelu_l131_40;
  wire                when_LeakyRelu_l133_40;
  wire                when_LeakyRelu_l131_41;
  wire                when_LeakyRelu_l133_41;
  wire                when_LeakyRelu_l131_42;
  wire                when_LeakyRelu_l133_42;
  wire                when_LeakyRelu_l131_43;
  wire                when_LeakyRelu_l133_43;
  wire                when_LeakyRelu_l131_44;
  wire                when_LeakyRelu_l133_44;
  wire                when_LeakyRelu_l131_45;
  wire                when_LeakyRelu_l133_45;
  wire                when_LeakyRelu_l131_46;
  wire                when_LeakyRelu_l133_46;
  wire                when_LeakyRelu_l131_47;
  wire                when_LeakyRelu_l133_47;
  wire       [15:0]   _zz_dataOut_2_1;
  wire                when_LeakyRelu_l155_2;
  wire                when_LeakyRelu_l157_2;
  reg        [7:0]    _zz_dataOut_3;
  reg        [15:0]   _zz_A_12;
  wire       [15:0]   _zz_when_LeakyRelu_l100_12;
  wire       [31:0]   _zz_when_LeakyRelu_l101_6;
  wire       [3:0]    _zz_when_LeakyRelu_l101_7;
  wire       [14:0]   _zz_A_13;
  wire       [14:0]   _zz_A_14;
  reg        [15:0]   _zz_when_LeakyRelu_l100_13;
  reg        [15:0]   _zz_when_LeakyRelu_l100_14;
  reg        [15:0]   _zz_when_LeakyRelu_l100_15;
  wire                when_LeakyRelu_l100_3;
  wire                when_LeakyRelu_l101_3;
  wire                when_LeakyRelu_l104_3;
  wire                when_LeakyRelu_l110_3;
  wire                when_LeakyRelu_l103_3;
  reg        [15:0]   _zz_A_15;
  reg        [15:0]   _zz_when_LeakyRelu_l100_15_regNext;
  wire                when_LeakyRelu_l127_3;
  wire                when_LeakyRelu_l131_48;
  wire                when_LeakyRelu_l133_48;
  wire                when_LeakyRelu_l131_49;
  wire                when_LeakyRelu_l133_49;
  wire                when_LeakyRelu_l131_50;
  wire                when_LeakyRelu_l133_50;
  wire                when_LeakyRelu_l131_51;
  wire                when_LeakyRelu_l133_51;
  wire                when_LeakyRelu_l131_52;
  wire                when_LeakyRelu_l133_52;
  wire                when_LeakyRelu_l131_53;
  wire                when_LeakyRelu_l133_53;
  wire                when_LeakyRelu_l131_54;
  wire                when_LeakyRelu_l133_54;
  wire                when_LeakyRelu_l131_55;
  wire                when_LeakyRelu_l133_55;
  wire                when_LeakyRelu_l131_56;
  wire                when_LeakyRelu_l133_56;
  wire                when_LeakyRelu_l131_57;
  wire                when_LeakyRelu_l133_57;
  wire                when_LeakyRelu_l131_58;
  wire                when_LeakyRelu_l133_58;
  wire                when_LeakyRelu_l131_59;
  wire                when_LeakyRelu_l133_59;
  wire                when_LeakyRelu_l131_60;
  wire                when_LeakyRelu_l133_60;
  wire                when_LeakyRelu_l131_61;
  wire                when_LeakyRelu_l133_61;
  wire                when_LeakyRelu_l131_62;
  wire                when_LeakyRelu_l133_62;
  wire                when_LeakyRelu_l131_63;
  wire                when_LeakyRelu_l133_63;
  wire       [15:0]   _zz_dataOut_3_1;
  wire                when_LeakyRelu_l155_3;
  wire                when_LeakyRelu_l157_3;
  reg        [7:0]    _zz_dataOut_4;
  reg        [15:0]   _zz_A_16;
  wire       [15:0]   _zz_when_LeakyRelu_l100_16;
  wire       [31:0]   _zz_when_LeakyRelu_l101_8;
  wire       [3:0]    _zz_when_LeakyRelu_l101_9;
  wire       [14:0]   _zz_A_17;
  wire       [14:0]   _zz_A_18;
  reg        [15:0]   _zz_when_LeakyRelu_l100_17;
  reg        [15:0]   _zz_when_LeakyRelu_l100_18;
  reg        [15:0]   _zz_when_LeakyRelu_l100_19;
  wire                when_LeakyRelu_l100_4;
  wire                when_LeakyRelu_l101_4;
  wire                when_LeakyRelu_l104_4;
  wire                when_LeakyRelu_l110_4;
  wire                when_LeakyRelu_l103_4;
  reg        [15:0]   _zz_A_19;
  reg        [15:0]   _zz_when_LeakyRelu_l100_19_regNext;
  wire                when_LeakyRelu_l127_4;
  wire                when_LeakyRelu_l131_64;
  wire                when_LeakyRelu_l133_64;
  wire                when_LeakyRelu_l131_65;
  wire                when_LeakyRelu_l133_65;
  wire                when_LeakyRelu_l131_66;
  wire                when_LeakyRelu_l133_66;
  wire                when_LeakyRelu_l131_67;
  wire                when_LeakyRelu_l133_67;
  wire                when_LeakyRelu_l131_68;
  wire                when_LeakyRelu_l133_68;
  wire                when_LeakyRelu_l131_69;
  wire                when_LeakyRelu_l133_69;
  wire                when_LeakyRelu_l131_70;
  wire                when_LeakyRelu_l133_70;
  wire                when_LeakyRelu_l131_71;
  wire                when_LeakyRelu_l133_71;
  wire                when_LeakyRelu_l131_72;
  wire                when_LeakyRelu_l133_72;
  wire                when_LeakyRelu_l131_73;
  wire                when_LeakyRelu_l133_73;
  wire                when_LeakyRelu_l131_74;
  wire                when_LeakyRelu_l133_74;
  wire                when_LeakyRelu_l131_75;
  wire                when_LeakyRelu_l133_75;
  wire                when_LeakyRelu_l131_76;
  wire                when_LeakyRelu_l133_76;
  wire                when_LeakyRelu_l131_77;
  wire                when_LeakyRelu_l133_77;
  wire                when_LeakyRelu_l131_78;
  wire                when_LeakyRelu_l133_78;
  wire                when_LeakyRelu_l131_79;
  wire                when_LeakyRelu_l133_79;
  wire       [15:0]   _zz_dataOut_4_1;
  wire                when_LeakyRelu_l155_4;
  wire                when_LeakyRelu_l157_4;
  reg        [7:0]    _zz_dataOut_5;
  reg        [15:0]   _zz_A_20;
  wire       [15:0]   _zz_when_LeakyRelu_l100_20;
  wire       [31:0]   _zz_when_LeakyRelu_l101_10;
  wire       [3:0]    _zz_when_LeakyRelu_l101_11;
  wire       [14:0]   _zz_A_21;
  wire       [14:0]   _zz_A_22;
  reg        [15:0]   _zz_when_LeakyRelu_l100_21;
  reg        [15:0]   _zz_when_LeakyRelu_l100_22;
  reg        [15:0]   _zz_when_LeakyRelu_l100_23;
  wire                when_LeakyRelu_l100_5;
  wire                when_LeakyRelu_l101_5;
  wire                when_LeakyRelu_l104_5;
  wire                when_LeakyRelu_l110_5;
  wire                when_LeakyRelu_l103_5;
  reg        [15:0]   _zz_A_23;
  reg        [15:0]   _zz_when_LeakyRelu_l100_23_regNext;
  wire                when_LeakyRelu_l127_5;
  wire                when_LeakyRelu_l131_80;
  wire                when_LeakyRelu_l133_80;
  wire                when_LeakyRelu_l131_81;
  wire                when_LeakyRelu_l133_81;
  wire                when_LeakyRelu_l131_82;
  wire                when_LeakyRelu_l133_82;
  wire                when_LeakyRelu_l131_83;
  wire                when_LeakyRelu_l133_83;
  wire                when_LeakyRelu_l131_84;
  wire                when_LeakyRelu_l133_84;
  wire                when_LeakyRelu_l131_85;
  wire                when_LeakyRelu_l133_85;
  wire                when_LeakyRelu_l131_86;
  wire                when_LeakyRelu_l133_86;
  wire                when_LeakyRelu_l131_87;
  wire                when_LeakyRelu_l133_87;
  wire                when_LeakyRelu_l131_88;
  wire                when_LeakyRelu_l133_88;
  wire                when_LeakyRelu_l131_89;
  wire                when_LeakyRelu_l133_89;
  wire                when_LeakyRelu_l131_90;
  wire                when_LeakyRelu_l133_90;
  wire                when_LeakyRelu_l131_91;
  wire                when_LeakyRelu_l133_91;
  wire                when_LeakyRelu_l131_92;
  wire                when_LeakyRelu_l133_92;
  wire                when_LeakyRelu_l131_93;
  wire                when_LeakyRelu_l133_93;
  wire                when_LeakyRelu_l131_94;
  wire                when_LeakyRelu_l133_94;
  wire                when_LeakyRelu_l131_95;
  wire                when_LeakyRelu_l133_95;
  wire       [15:0]   _zz_dataOut_5_1;
  wire                when_LeakyRelu_l155_5;
  wire                when_LeakyRelu_l157_5;
  reg        [7:0]    _zz_dataOut_6;
  reg        [15:0]   _zz_A_24;
  wire       [15:0]   _zz_when_LeakyRelu_l100_24;
  wire       [31:0]   _zz_when_LeakyRelu_l101_12;
  wire       [3:0]    _zz_when_LeakyRelu_l101_13;
  wire       [14:0]   _zz_A_25;
  wire       [14:0]   _zz_A_26;
  reg        [15:0]   _zz_when_LeakyRelu_l100_25;
  reg        [15:0]   _zz_when_LeakyRelu_l100_26;
  reg        [15:0]   _zz_when_LeakyRelu_l100_27;
  wire                when_LeakyRelu_l100_6;
  wire                when_LeakyRelu_l101_6;
  wire                when_LeakyRelu_l104_6;
  wire                when_LeakyRelu_l110_6;
  wire                when_LeakyRelu_l103_6;
  reg        [15:0]   _zz_A_27;
  reg        [15:0]   _zz_when_LeakyRelu_l100_27_regNext;
  wire                when_LeakyRelu_l127_6;
  wire                when_LeakyRelu_l131_96;
  wire                when_LeakyRelu_l133_96;
  wire                when_LeakyRelu_l131_97;
  wire                when_LeakyRelu_l133_97;
  wire                when_LeakyRelu_l131_98;
  wire                when_LeakyRelu_l133_98;
  wire                when_LeakyRelu_l131_99;
  wire                when_LeakyRelu_l133_99;
  wire                when_LeakyRelu_l131_100;
  wire                when_LeakyRelu_l133_100;
  wire                when_LeakyRelu_l131_101;
  wire                when_LeakyRelu_l133_101;
  wire                when_LeakyRelu_l131_102;
  wire                when_LeakyRelu_l133_102;
  wire                when_LeakyRelu_l131_103;
  wire                when_LeakyRelu_l133_103;
  wire                when_LeakyRelu_l131_104;
  wire                when_LeakyRelu_l133_104;
  wire                when_LeakyRelu_l131_105;
  wire                when_LeakyRelu_l133_105;
  wire                when_LeakyRelu_l131_106;
  wire                when_LeakyRelu_l133_106;
  wire                when_LeakyRelu_l131_107;
  wire                when_LeakyRelu_l133_107;
  wire                when_LeakyRelu_l131_108;
  wire                when_LeakyRelu_l133_108;
  wire                when_LeakyRelu_l131_109;
  wire                when_LeakyRelu_l133_109;
  wire                when_LeakyRelu_l131_110;
  wire                when_LeakyRelu_l133_110;
  wire                when_LeakyRelu_l131_111;
  wire                when_LeakyRelu_l133_111;
  wire       [15:0]   _zz_dataOut_6_1;
  wire                when_LeakyRelu_l155_6;
  wire                when_LeakyRelu_l157_6;
  reg        [7:0]    _zz_dataOut_7;
  reg        [15:0]   _zz_A_28;
  wire       [15:0]   _zz_when_LeakyRelu_l100_28;
  wire       [31:0]   _zz_when_LeakyRelu_l101_14;
  wire       [3:0]    _zz_when_LeakyRelu_l101_15;
  wire       [14:0]   _zz_A_29;
  wire       [14:0]   _zz_A_30;
  reg        [15:0]   _zz_when_LeakyRelu_l100_29;
  reg        [15:0]   _zz_when_LeakyRelu_l100_30;
  reg        [15:0]   _zz_when_LeakyRelu_l100_31;
  wire                when_LeakyRelu_l100_7;
  wire                when_LeakyRelu_l101_7;
  wire                when_LeakyRelu_l104_7;
  wire                when_LeakyRelu_l110_7;
  wire                when_LeakyRelu_l103_7;
  reg        [15:0]   _zz_A_31;
  reg        [15:0]   _zz_when_LeakyRelu_l100_31_regNext;
  wire                when_LeakyRelu_l127_7;
  wire                when_LeakyRelu_l131_112;
  wire                when_LeakyRelu_l133_112;
  wire                when_LeakyRelu_l131_113;
  wire                when_LeakyRelu_l133_113;
  wire                when_LeakyRelu_l131_114;
  wire                when_LeakyRelu_l133_114;
  wire                when_LeakyRelu_l131_115;
  wire                when_LeakyRelu_l133_115;
  wire                when_LeakyRelu_l131_116;
  wire                when_LeakyRelu_l133_116;
  wire                when_LeakyRelu_l131_117;
  wire                when_LeakyRelu_l133_117;
  wire                when_LeakyRelu_l131_118;
  wire                when_LeakyRelu_l133_118;
  wire                when_LeakyRelu_l131_119;
  wire                when_LeakyRelu_l133_119;
  wire                when_LeakyRelu_l131_120;
  wire                when_LeakyRelu_l133_120;
  wire                when_LeakyRelu_l131_121;
  wire                when_LeakyRelu_l133_121;
  wire                when_LeakyRelu_l131_122;
  wire                when_LeakyRelu_l133_122;
  wire                when_LeakyRelu_l131_123;
  wire                when_LeakyRelu_l133_123;
  wire                when_LeakyRelu_l131_124;
  wire                when_LeakyRelu_l133_124;
  wire                when_LeakyRelu_l131_125;
  wire                when_LeakyRelu_l133_125;
  wire                when_LeakyRelu_l131_126;
  wire                when_LeakyRelu_l133_126;
  wire                when_LeakyRelu_l131_127;
  wire                when_LeakyRelu_l133_127;
  wire       [15:0]   _zz_dataOut_7_1;
  wire                when_LeakyRelu_l155_7;
  wire                when_LeakyRelu_l157_7;
  reg        [7:0]    _zz_dataOut_8;
  reg        [15:0]   _zz_A_32;
  wire       [15:0]   _zz_when_LeakyRelu_l100_32;
  wire       [31:0]   _zz_when_LeakyRelu_l101_16;
  wire       [3:0]    _zz_when_LeakyRelu_l101_17;
  wire       [14:0]   _zz_A_33;
  wire       [14:0]   _zz_A_34;
  reg        [15:0]   _zz_when_LeakyRelu_l100_33;
  reg        [15:0]   _zz_when_LeakyRelu_l100_34;
  reg        [15:0]   _zz_when_LeakyRelu_l100_35;
  wire                when_LeakyRelu_l100_8;
  wire                when_LeakyRelu_l101_8;
  wire                when_LeakyRelu_l104_8;
  wire                when_LeakyRelu_l110_8;
  wire                when_LeakyRelu_l103_8;
  reg        [15:0]   _zz_A_35;
  reg        [15:0]   _zz_when_LeakyRelu_l100_35_regNext;
  wire                when_LeakyRelu_l127_8;
  wire                when_LeakyRelu_l131_128;
  wire                when_LeakyRelu_l133_128;
  wire                when_LeakyRelu_l131_129;
  wire                when_LeakyRelu_l133_129;
  wire                when_LeakyRelu_l131_130;
  wire                when_LeakyRelu_l133_130;
  wire                when_LeakyRelu_l131_131;
  wire                when_LeakyRelu_l133_131;
  wire                when_LeakyRelu_l131_132;
  wire                when_LeakyRelu_l133_132;
  wire                when_LeakyRelu_l131_133;
  wire                when_LeakyRelu_l133_133;
  wire                when_LeakyRelu_l131_134;
  wire                when_LeakyRelu_l133_134;
  wire                when_LeakyRelu_l131_135;
  wire                when_LeakyRelu_l133_135;
  wire                when_LeakyRelu_l131_136;
  wire                when_LeakyRelu_l133_136;
  wire                when_LeakyRelu_l131_137;
  wire                when_LeakyRelu_l133_137;
  wire                when_LeakyRelu_l131_138;
  wire                when_LeakyRelu_l133_138;
  wire                when_LeakyRelu_l131_139;
  wire                when_LeakyRelu_l133_139;
  wire                when_LeakyRelu_l131_140;
  wire                when_LeakyRelu_l133_140;
  wire                when_LeakyRelu_l131_141;
  wire                when_LeakyRelu_l133_141;
  wire                when_LeakyRelu_l131_142;
  wire                when_LeakyRelu_l133_142;
  wire                when_LeakyRelu_l131_143;
  wire                when_LeakyRelu_l133_143;
  wire       [15:0]   _zz_dataOut_8_1;
  wire                when_LeakyRelu_l155_8;
  wire                when_LeakyRelu_l157_8;
  reg        [7:0]    _zz_dataOut_9;
  reg        [15:0]   _zz_A_36;
  wire       [15:0]   _zz_when_LeakyRelu_l100_36;
  wire       [31:0]   _zz_when_LeakyRelu_l101_18;
  wire       [3:0]    _zz_when_LeakyRelu_l101_19;
  wire       [14:0]   _zz_A_37;
  wire       [14:0]   _zz_A_38;
  reg        [15:0]   _zz_when_LeakyRelu_l100_37;
  reg        [15:0]   _zz_when_LeakyRelu_l100_38;
  reg        [15:0]   _zz_when_LeakyRelu_l100_39;
  wire                when_LeakyRelu_l100_9;
  wire                when_LeakyRelu_l101_9;
  wire                when_LeakyRelu_l104_9;
  wire                when_LeakyRelu_l110_9;
  wire                when_LeakyRelu_l103_9;
  reg        [15:0]   _zz_A_39;
  reg        [15:0]   _zz_when_LeakyRelu_l100_39_regNext;
  wire                when_LeakyRelu_l127_9;
  wire                when_LeakyRelu_l131_144;
  wire                when_LeakyRelu_l133_144;
  wire                when_LeakyRelu_l131_145;
  wire                when_LeakyRelu_l133_145;
  wire                when_LeakyRelu_l131_146;
  wire                when_LeakyRelu_l133_146;
  wire                when_LeakyRelu_l131_147;
  wire                when_LeakyRelu_l133_147;
  wire                when_LeakyRelu_l131_148;
  wire                when_LeakyRelu_l133_148;
  wire                when_LeakyRelu_l131_149;
  wire                when_LeakyRelu_l133_149;
  wire                when_LeakyRelu_l131_150;
  wire                when_LeakyRelu_l133_150;
  wire                when_LeakyRelu_l131_151;
  wire                when_LeakyRelu_l133_151;
  wire                when_LeakyRelu_l131_152;
  wire                when_LeakyRelu_l133_152;
  wire                when_LeakyRelu_l131_153;
  wire                when_LeakyRelu_l133_153;
  wire                when_LeakyRelu_l131_154;
  wire                when_LeakyRelu_l133_154;
  wire                when_LeakyRelu_l131_155;
  wire                when_LeakyRelu_l133_155;
  wire                when_LeakyRelu_l131_156;
  wire                when_LeakyRelu_l133_156;
  wire                when_LeakyRelu_l131_157;
  wire                when_LeakyRelu_l133_157;
  wire                when_LeakyRelu_l131_158;
  wire                when_LeakyRelu_l133_158;
  wire                when_LeakyRelu_l131_159;
  wire                when_LeakyRelu_l133_159;
  wire       [15:0]   _zz_dataOut_9_1;
  wire                when_LeakyRelu_l155_9;
  wire                when_LeakyRelu_l157_9;
  reg        [7:0]    _zz_dataOut_10;
  reg        [15:0]   _zz_A_40;
  wire       [15:0]   _zz_when_LeakyRelu_l100_40;
  wire       [31:0]   _zz_when_LeakyRelu_l101_20;
  wire       [3:0]    _zz_when_LeakyRelu_l101_21;
  wire       [14:0]   _zz_A_41;
  wire       [14:0]   _zz_A_42;
  reg        [15:0]   _zz_when_LeakyRelu_l100_41;
  reg        [15:0]   _zz_when_LeakyRelu_l100_42;
  reg        [15:0]   _zz_when_LeakyRelu_l100_43;
  wire                when_LeakyRelu_l100_10;
  wire                when_LeakyRelu_l101_10;
  wire                when_LeakyRelu_l104_10;
  wire                when_LeakyRelu_l110_10;
  wire                when_LeakyRelu_l103_10;
  reg        [15:0]   _zz_A_43;
  reg        [15:0]   _zz_when_LeakyRelu_l100_43_regNext;
  wire                when_LeakyRelu_l127_10;
  wire                when_LeakyRelu_l131_160;
  wire                when_LeakyRelu_l133_160;
  wire                when_LeakyRelu_l131_161;
  wire                when_LeakyRelu_l133_161;
  wire                when_LeakyRelu_l131_162;
  wire                when_LeakyRelu_l133_162;
  wire                when_LeakyRelu_l131_163;
  wire                when_LeakyRelu_l133_163;
  wire                when_LeakyRelu_l131_164;
  wire                when_LeakyRelu_l133_164;
  wire                when_LeakyRelu_l131_165;
  wire                when_LeakyRelu_l133_165;
  wire                when_LeakyRelu_l131_166;
  wire                when_LeakyRelu_l133_166;
  wire                when_LeakyRelu_l131_167;
  wire                when_LeakyRelu_l133_167;
  wire                when_LeakyRelu_l131_168;
  wire                when_LeakyRelu_l133_168;
  wire                when_LeakyRelu_l131_169;
  wire                when_LeakyRelu_l133_169;
  wire                when_LeakyRelu_l131_170;
  wire                when_LeakyRelu_l133_170;
  wire                when_LeakyRelu_l131_171;
  wire                when_LeakyRelu_l133_171;
  wire                when_LeakyRelu_l131_172;
  wire                when_LeakyRelu_l133_172;
  wire                when_LeakyRelu_l131_173;
  wire                when_LeakyRelu_l133_173;
  wire                when_LeakyRelu_l131_174;
  wire                when_LeakyRelu_l133_174;
  wire                when_LeakyRelu_l131_175;
  wire                when_LeakyRelu_l133_175;
  wire       [15:0]   _zz_dataOut_10_1;
  wire                when_LeakyRelu_l155_10;
  wire                when_LeakyRelu_l157_10;
  reg        [7:0]    _zz_dataOut_11;
  reg        [15:0]   _zz_A_44;
  wire       [15:0]   _zz_when_LeakyRelu_l100_44;
  wire       [31:0]   _zz_when_LeakyRelu_l101_22;
  wire       [3:0]    _zz_when_LeakyRelu_l101_23;
  wire       [14:0]   _zz_A_45;
  wire       [14:0]   _zz_A_46;
  reg        [15:0]   _zz_when_LeakyRelu_l100_45;
  reg        [15:0]   _zz_when_LeakyRelu_l100_46;
  reg        [15:0]   _zz_when_LeakyRelu_l100_47;
  wire                when_LeakyRelu_l100_11;
  wire                when_LeakyRelu_l101_11;
  wire                when_LeakyRelu_l104_11;
  wire                when_LeakyRelu_l110_11;
  wire                when_LeakyRelu_l103_11;
  reg        [15:0]   _zz_A_47;
  reg        [15:0]   _zz_when_LeakyRelu_l100_47_regNext;
  wire                when_LeakyRelu_l127_11;
  wire                when_LeakyRelu_l131_176;
  wire                when_LeakyRelu_l133_176;
  wire                when_LeakyRelu_l131_177;
  wire                when_LeakyRelu_l133_177;
  wire                when_LeakyRelu_l131_178;
  wire                when_LeakyRelu_l133_178;
  wire                when_LeakyRelu_l131_179;
  wire                when_LeakyRelu_l133_179;
  wire                when_LeakyRelu_l131_180;
  wire                when_LeakyRelu_l133_180;
  wire                when_LeakyRelu_l131_181;
  wire                when_LeakyRelu_l133_181;
  wire                when_LeakyRelu_l131_182;
  wire                when_LeakyRelu_l133_182;
  wire                when_LeakyRelu_l131_183;
  wire                when_LeakyRelu_l133_183;
  wire                when_LeakyRelu_l131_184;
  wire                when_LeakyRelu_l133_184;
  wire                when_LeakyRelu_l131_185;
  wire                when_LeakyRelu_l133_185;
  wire                when_LeakyRelu_l131_186;
  wire                when_LeakyRelu_l133_186;
  wire                when_LeakyRelu_l131_187;
  wire                when_LeakyRelu_l133_187;
  wire                when_LeakyRelu_l131_188;
  wire                when_LeakyRelu_l133_188;
  wire                when_LeakyRelu_l131_189;
  wire                when_LeakyRelu_l133_189;
  wire                when_LeakyRelu_l131_190;
  wire                when_LeakyRelu_l133_190;
  wire                when_LeakyRelu_l131_191;
  wire                when_LeakyRelu_l133_191;
  wire       [15:0]   _zz_dataOut_11_1;
  wire                when_LeakyRelu_l155_11;
  wire                when_LeakyRelu_l157_11;
  reg        [7:0]    _zz_dataOut_12;
  reg        [15:0]   _zz_A_48;
  wire       [15:0]   _zz_when_LeakyRelu_l100_48;
  wire       [31:0]   _zz_when_LeakyRelu_l101_24;
  wire       [3:0]    _zz_when_LeakyRelu_l101_25;
  wire       [14:0]   _zz_A_49;
  wire       [14:0]   _zz_A_50;
  reg        [15:0]   _zz_when_LeakyRelu_l100_49;
  reg        [15:0]   _zz_when_LeakyRelu_l100_50;
  reg        [15:0]   _zz_when_LeakyRelu_l100_51;
  wire                when_LeakyRelu_l100_12;
  wire                when_LeakyRelu_l101_12;
  wire                when_LeakyRelu_l104_12;
  wire                when_LeakyRelu_l110_12;
  wire                when_LeakyRelu_l103_12;
  reg        [15:0]   _zz_A_51;
  reg        [15:0]   _zz_when_LeakyRelu_l100_51_regNext;
  wire                when_LeakyRelu_l127_12;
  wire                when_LeakyRelu_l131_192;
  wire                when_LeakyRelu_l133_192;
  wire                when_LeakyRelu_l131_193;
  wire                when_LeakyRelu_l133_193;
  wire                when_LeakyRelu_l131_194;
  wire                when_LeakyRelu_l133_194;
  wire                when_LeakyRelu_l131_195;
  wire                when_LeakyRelu_l133_195;
  wire                when_LeakyRelu_l131_196;
  wire                when_LeakyRelu_l133_196;
  wire                when_LeakyRelu_l131_197;
  wire                when_LeakyRelu_l133_197;
  wire                when_LeakyRelu_l131_198;
  wire                when_LeakyRelu_l133_198;
  wire                when_LeakyRelu_l131_199;
  wire                when_LeakyRelu_l133_199;
  wire                when_LeakyRelu_l131_200;
  wire                when_LeakyRelu_l133_200;
  wire                when_LeakyRelu_l131_201;
  wire                when_LeakyRelu_l133_201;
  wire                when_LeakyRelu_l131_202;
  wire                when_LeakyRelu_l133_202;
  wire                when_LeakyRelu_l131_203;
  wire                when_LeakyRelu_l133_203;
  wire                when_LeakyRelu_l131_204;
  wire                when_LeakyRelu_l133_204;
  wire                when_LeakyRelu_l131_205;
  wire                when_LeakyRelu_l133_205;
  wire                when_LeakyRelu_l131_206;
  wire                when_LeakyRelu_l133_206;
  wire                when_LeakyRelu_l131_207;
  wire                when_LeakyRelu_l133_207;
  wire       [15:0]   _zz_dataOut_12_1;
  wire                when_LeakyRelu_l155_12;
  wire                when_LeakyRelu_l157_12;
  reg        [7:0]    _zz_dataOut_13;
  reg        [15:0]   _zz_A_52;
  wire       [15:0]   _zz_when_LeakyRelu_l100_52;
  wire       [31:0]   _zz_when_LeakyRelu_l101_26;
  wire       [3:0]    _zz_when_LeakyRelu_l101_27;
  wire       [14:0]   _zz_A_53;
  wire       [14:0]   _zz_A_54;
  reg        [15:0]   _zz_when_LeakyRelu_l100_53;
  reg        [15:0]   _zz_when_LeakyRelu_l100_54;
  reg        [15:0]   _zz_when_LeakyRelu_l100_55;
  wire                when_LeakyRelu_l100_13;
  wire                when_LeakyRelu_l101_13;
  wire                when_LeakyRelu_l104_13;
  wire                when_LeakyRelu_l110_13;
  wire                when_LeakyRelu_l103_13;
  reg        [15:0]   _zz_A_55;
  reg        [15:0]   _zz_when_LeakyRelu_l100_55_regNext;
  wire                when_LeakyRelu_l127_13;
  wire                when_LeakyRelu_l131_208;
  wire                when_LeakyRelu_l133_208;
  wire                when_LeakyRelu_l131_209;
  wire                when_LeakyRelu_l133_209;
  wire                when_LeakyRelu_l131_210;
  wire                when_LeakyRelu_l133_210;
  wire                when_LeakyRelu_l131_211;
  wire                when_LeakyRelu_l133_211;
  wire                when_LeakyRelu_l131_212;
  wire                when_LeakyRelu_l133_212;
  wire                when_LeakyRelu_l131_213;
  wire                when_LeakyRelu_l133_213;
  wire                when_LeakyRelu_l131_214;
  wire                when_LeakyRelu_l133_214;
  wire                when_LeakyRelu_l131_215;
  wire                when_LeakyRelu_l133_215;
  wire                when_LeakyRelu_l131_216;
  wire                when_LeakyRelu_l133_216;
  wire                when_LeakyRelu_l131_217;
  wire                when_LeakyRelu_l133_217;
  wire                when_LeakyRelu_l131_218;
  wire                when_LeakyRelu_l133_218;
  wire                when_LeakyRelu_l131_219;
  wire                when_LeakyRelu_l133_219;
  wire                when_LeakyRelu_l131_220;
  wire                when_LeakyRelu_l133_220;
  wire                when_LeakyRelu_l131_221;
  wire                when_LeakyRelu_l133_221;
  wire                when_LeakyRelu_l131_222;
  wire                when_LeakyRelu_l133_222;
  wire                when_LeakyRelu_l131_223;
  wire                when_LeakyRelu_l133_223;
  wire       [15:0]   _zz_dataOut_13_1;
  wire                when_LeakyRelu_l155_13;
  wire                when_LeakyRelu_l157_13;
  reg        [7:0]    _zz_dataOut_14;
  reg        [15:0]   _zz_A_56;
  wire       [15:0]   _zz_when_LeakyRelu_l100_56;
  wire       [31:0]   _zz_when_LeakyRelu_l101_28;
  wire       [3:0]    _zz_when_LeakyRelu_l101_29;
  wire       [14:0]   _zz_A_57;
  wire       [14:0]   _zz_A_58;
  reg        [15:0]   _zz_when_LeakyRelu_l100_57;
  reg        [15:0]   _zz_when_LeakyRelu_l100_58;
  reg        [15:0]   _zz_when_LeakyRelu_l100_59;
  wire                when_LeakyRelu_l100_14;
  wire                when_LeakyRelu_l101_14;
  wire                when_LeakyRelu_l104_14;
  wire                when_LeakyRelu_l110_14;
  wire                when_LeakyRelu_l103_14;
  reg        [15:0]   _zz_A_59;
  reg        [15:0]   _zz_when_LeakyRelu_l100_59_regNext;
  wire                when_LeakyRelu_l127_14;
  wire                when_LeakyRelu_l131_224;
  wire                when_LeakyRelu_l133_224;
  wire                when_LeakyRelu_l131_225;
  wire                when_LeakyRelu_l133_225;
  wire                when_LeakyRelu_l131_226;
  wire                when_LeakyRelu_l133_226;
  wire                when_LeakyRelu_l131_227;
  wire                when_LeakyRelu_l133_227;
  wire                when_LeakyRelu_l131_228;
  wire                when_LeakyRelu_l133_228;
  wire                when_LeakyRelu_l131_229;
  wire                when_LeakyRelu_l133_229;
  wire                when_LeakyRelu_l131_230;
  wire                when_LeakyRelu_l133_230;
  wire                when_LeakyRelu_l131_231;
  wire                when_LeakyRelu_l133_231;
  wire                when_LeakyRelu_l131_232;
  wire                when_LeakyRelu_l133_232;
  wire                when_LeakyRelu_l131_233;
  wire                when_LeakyRelu_l133_233;
  wire                when_LeakyRelu_l131_234;
  wire                when_LeakyRelu_l133_234;
  wire                when_LeakyRelu_l131_235;
  wire                when_LeakyRelu_l133_235;
  wire                when_LeakyRelu_l131_236;
  wire                when_LeakyRelu_l133_236;
  wire                when_LeakyRelu_l131_237;
  wire                when_LeakyRelu_l133_237;
  wire                when_LeakyRelu_l131_238;
  wire                when_LeakyRelu_l133_238;
  wire                when_LeakyRelu_l131_239;
  wire                when_LeakyRelu_l133_239;
  wire       [15:0]   _zz_dataOut_14_1;
  wire                when_LeakyRelu_l155_14;
  wire                when_LeakyRelu_l157_14;
  reg        [7:0]    _zz_dataOut_15;
  reg        [15:0]   _zz_A_60;
  wire       [15:0]   _zz_when_LeakyRelu_l100_60;
  wire       [31:0]   _zz_when_LeakyRelu_l101_30;
  wire       [3:0]    _zz_when_LeakyRelu_l101_31;
  wire       [14:0]   _zz_A_61;
  wire       [14:0]   _zz_A_62;
  reg        [15:0]   _zz_when_LeakyRelu_l100_61;
  reg        [15:0]   _zz_when_LeakyRelu_l100_62;
  reg        [15:0]   _zz_when_LeakyRelu_l100_63;
  wire                when_LeakyRelu_l100_15;
  wire                when_LeakyRelu_l101_15;
  wire                when_LeakyRelu_l104_15;
  wire                when_LeakyRelu_l110_15;
  wire                when_LeakyRelu_l103_15;
  reg        [15:0]   _zz_A_63;
  reg        [15:0]   _zz_when_LeakyRelu_l100_63_regNext;
  wire                when_LeakyRelu_l127_15;
  wire                when_LeakyRelu_l131_240;
  wire                when_LeakyRelu_l133_240;
  wire                when_LeakyRelu_l131_241;
  wire                when_LeakyRelu_l133_241;
  wire                when_LeakyRelu_l131_242;
  wire                when_LeakyRelu_l133_242;
  wire                when_LeakyRelu_l131_243;
  wire                when_LeakyRelu_l133_243;
  wire                when_LeakyRelu_l131_244;
  wire                when_LeakyRelu_l133_244;
  wire                when_LeakyRelu_l131_245;
  wire                when_LeakyRelu_l133_245;
  wire                when_LeakyRelu_l131_246;
  wire                when_LeakyRelu_l133_246;
  wire                when_LeakyRelu_l131_247;
  wire                when_LeakyRelu_l133_247;
  wire                when_LeakyRelu_l131_248;
  wire                when_LeakyRelu_l133_248;
  wire                when_LeakyRelu_l131_249;
  wire                when_LeakyRelu_l133_249;
  wire                when_LeakyRelu_l131_250;
  wire                when_LeakyRelu_l133_250;
  wire                when_LeakyRelu_l131_251;
  wire                when_LeakyRelu_l133_251;
  wire                when_LeakyRelu_l131_252;
  wire                when_LeakyRelu_l133_252;
  wire                when_LeakyRelu_l131_253;
  wire                when_LeakyRelu_l133_253;
  wire                when_LeakyRelu_l131_254;
  wire                when_LeakyRelu_l133_254;
  wire                when_LeakyRelu_l131_255;
  wire                when_LeakyRelu_l133_255;
  wire       [15:0]   _zz_dataOut_15_1;
  wire                when_LeakyRelu_l155_15;
  wire                when_LeakyRelu_l157_15;

  assign _zz__zz_A_1 = (_zz_when_LeakyRelu_l101 >>> 17);
  assign _zz__zz_A_1_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_32 = 4'b0000;
  assign _zz_1 = 16'hfffb;
  assign _zz_2 = 16'hfff1;
  assign _zz_3 = 16'hffe7;
  assign _zz_4 = 16'hffdd;
  assign _zz_5 = 16'hffd3;
  assign _zz_6 = 16'hffc9;
  assign _zz_7 = 16'hffbf;
  assign _zz_8 = 16'hffb5;
  assign _zz_9 = 16'hffab;
  assign _zz_10 = 16'hffa1;
  assign _zz_11 = 16'hff97;
  assign _zz_12 = 16'hff8d;
  assign _zz_13 = 16'hff83;
  assign _zz_14 = 16'hff79;
  assign _zz_15 = 16'hff6f;
  assign _zz_16 = 16'hff65;
  assign _zz__zz_A_3 = 16'h0001;
  assign _zz__zz_A_3_1 = 16'h0001;
  assign _zz__zz_A_3_2 = 16'h0001;
  assign _zz__zz_A_3_3 = 16'h0001;
  assign _zz__zz_A_3_4 = 16'h0001;
  assign _zz__zz_A_3_5 = 16'h0001;
  assign _zz__zz_A_3_6 = 16'h0001;
  assign _zz__zz_A_3_7 = 16'h0001;
  assign _zz__zz_A_3_8 = 16'h0001;
  assign _zz__zz_A_3_9 = 16'h0001;
  assign _zz__zz_A_3_10 = 16'h0001;
  assign _zz__zz_A_3_11 = 16'h0001;
  assign _zz__zz_A_3_12 = 16'h0001;
  assign _zz__zz_A_3_13 = 16'h0001;
  assign _zz__zz_A_3_14 = 16'h0001;
  assign _zz__zz_A_3_15 = 16'h0001;
  assign _zz__zz_A_3_16 = 16'h0001;
  assign _zz__zz_A_3_17 = 16'h0001;
  assign _zz__zz_A_3_18 = 16'h0001;
  assign _zz__zz_A_3_19 = 16'h0001;
  assign _zz__zz_A_3_20 = 16'h0001;
  assign _zz__zz_A_3_21 = 16'h0001;
  assign _zz__zz_A_3_22 = 16'h0001;
  assign _zz__zz_A_3_23 = 16'h0001;
  assign _zz__zz_A_3_24 = 16'h0001;
  assign _zz__zz_A_3_25 = 16'h0001;
  assign _zz__zz_A_3_26 = 16'h0001;
  assign _zz__zz_A_3_27 = 16'h0001;
  assign _zz__zz_A_3_28 = 16'h0001;
  assign _zz__zz_A_3_29 = 16'h0001;
  assign _zz__zz_A_3_30 = 16'h0001;
  assign _zz__zz_A_3_31 = 16'h0001;
  assign _zz__zz_dataOut_0 = _zz_dataOut_0_1;
  assign _zz_when_LeakyRelu_l157 = 16'h00ff;
  assign _zz__zz_A_5 = (_zz_when_LeakyRelu_l101_2 >>> 17);
  assign _zz__zz_A_5_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_1_1 = 4'b0000;
  assign _zz_17 = 16'hfffb;
  assign _zz_18 = 16'hfff1;
  assign _zz_19 = 16'hffe7;
  assign _zz_20 = 16'hffdd;
  assign _zz_21 = 16'hffd3;
  assign _zz_22 = 16'hffc9;
  assign _zz_23 = 16'hffbf;
  assign _zz_24 = 16'hffb5;
  assign _zz_25 = 16'hffab;
  assign _zz_26 = 16'hffa1;
  assign _zz_27 = 16'hff97;
  assign _zz_28 = 16'hff8d;
  assign _zz_29 = 16'hff83;
  assign _zz_30 = 16'hff79;
  assign _zz_31 = 16'hff6f;
  assign _zz_32 = 16'hff65;
  assign _zz__zz_A_7 = 16'h0001;
  assign _zz__zz_A_7_1 = 16'h0001;
  assign _zz__zz_A_7_2 = 16'h0001;
  assign _zz__zz_A_7_3 = 16'h0001;
  assign _zz__zz_A_7_4 = 16'h0001;
  assign _zz__zz_A_7_5 = 16'h0001;
  assign _zz__zz_A_7_6 = 16'h0001;
  assign _zz__zz_A_7_7 = 16'h0001;
  assign _zz__zz_A_7_8 = 16'h0001;
  assign _zz__zz_A_7_9 = 16'h0001;
  assign _zz__zz_A_7_10 = 16'h0001;
  assign _zz__zz_A_7_11 = 16'h0001;
  assign _zz__zz_A_7_12 = 16'h0001;
  assign _zz__zz_A_7_13 = 16'h0001;
  assign _zz__zz_A_7_14 = 16'h0001;
  assign _zz__zz_A_7_15 = 16'h0001;
  assign _zz__zz_A_7_16 = 16'h0001;
  assign _zz__zz_A_7_17 = 16'h0001;
  assign _zz__zz_A_7_18 = 16'h0001;
  assign _zz__zz_A_7_19 = 16'h0001;
  assign _zz__zz_A_7_20 = 16'h0001;
  assign _zz__zz_A_7_21 = 16'h0001;
  assign _zz__zz_A_7_22 = 16'h0001;
  assign _zz__zz_A_7_23 = 16'h0001;
  assign _zz__zz_A_7_24 = 16'h0001;
  assign _zz__zz_A_7_25 = 16'h0001;
  assign _zz__zz_A_7_26 = 16'h0001;
  assign _zz__zz_A_7_27 = 16'h0001;
  assign _zz__zz_A_7_28 = 16'h0001;
  assign _zz__zz_A_7_29 = 16'h0001;
  assign _zz__zz_A_7_30 = 16'h0001;
  assign _zz__zz_A_7_31 = 16'h0001;
  assign _zz__zz_dataOut_1 = _zz_dataOut_1_1;
  assign _zz_when_LeakyRelu_l157_1 = 16'h00ff;
  assign _zz__zz_A_9 = (_zz_when_LeakyRelu_l101_4 >>> 17);
  assign _zz__zz_A_9_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_2_1 = 4'b0000;
  assign _zz_33 = 16'hfffb;
  assign _zz_34 = 16'hfff1;
  assign _zz_35 = 16'hffe7;
  assign _zz_36 = 16'hffdd;
  assign _zz_37 = 16'hffd3;
  assign _zz_38 = 16'hffc9;
  assign _zz_39 = 16'hffbf;
  assign _zz_40 = 16'hffb5;
  assign _zz_41 = 16'hffab;
  assign _zz_42 = 16'hffa1;
  assign _zz_43 = 16'hff97;
  assign _zz_44 = 16'hff8d;
  assign _zz_45 = 16'hff83;
  assign _zz_46 = 16'hff79;
  assign _zz_47 = 16'hff6f;
  assign _zz_48 = 16'hff65;
  assign _zz__zz_A_11 = 16'h0001;
  assign _zz__zz_A_11_1 = 16'h0001;
  assign _zz__zz_A_11_2 = 16'h0001;
  assign _zz__zz_A_11_3 = 16'h0001;
  assign _zz__zz_A_11_4 = 16'h0001;
  assign _zz__zz_A_11_5 = 16'h0001;
  assign _zz__zz_A_11_6 = 16'h0001;
  assign _zz__zz_A_11_7 = 16'h0001;
  assign _zz__zz_A_11_8 = 16'h0001;
  assign _zz__zz_A_11_9 = 16'h0001;
  assign _zz__zz_A_11_10 = 16'h0001;
  assign _zz__zz_A_11_11 = 16'h0001;
  assign _zz__zz_A_11_12 = 16'h0001;
  assign _zz__zz_A_11_13 = 16'h0001;
  assign _zz__zz_A_11_14 = 16'h0001;
  assign _zz__zz_A_11_15 = 16'h0001;
  assign _zz__zz_A_11_16 = 16'h0001;
  assign _zz__zz_A_11_17 = 16'h0001;
  assign _zz__zz_A_11_18 = 16'h0001;
  assign _zz__zz_A_11_19 = 16'h0001;
  assign _zz__zz_A_11_20 = 16'h0001;
  assign _zz__zz_A_11_21 = 16'h0001;
  assign _zz__zz_A_11_22 = 16'h0001;
  assign _zz__zz_A_11_23 = 16'h0001;
  assign _zz__zz_A_11_24 = 16'h0001;
  assign _zz__zz_A_11_25 = 16'h0001;
  assign _zz__zz_A_11_26 = 16'h0001;
  assign _zz__zz_A_11_27 = 16'h0001;
  assign _zz__zz_A_11_28 = 16'h0001;
  assign _zz__zz_A_11_29 = 16'h0001;
  assign _zz__zz_A_11_30 = 16'h0001;
  assign _zz__zz_A_11_31 = 16'h0001;
  assign _zz__zz_dataOut_2 = _zz_dataOut_2_1;
  assign _zz_when_LeakyRelu_l157_2 = 16'h00ff;
  assign _zz__zz_A_13 = (_zz_when_LeakyRelu_l101_6 >>> 17);
  assign _zz__zz_A_13_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_3_1 = 4'b0000;
  assign _zz_49 = 16'hfffb;
  assign _zz_50 = 16'hfff1;
  assign _zz_51 = 16'hffe7;
  assign _zz_52 = 16'hffdd;
  assign _zz_53 = 16'hffd3;
  assign _zz_54 = 16'hffc9;
  assign _zz_55 = 16'hffbf;
  assign _zz_56 = 16'hffb5;
  assign _zz_57 = 16'hffab;
  assign _zz_58 = 16'hffa1;
  assign _zz_59 = 16'hff97;
  assign _zz_60 = 16'hff8d;
  assign _zz_61 = 16'hff83;
  assign _zz_62 = 16'hff79;
  assign _zz_63 = 16'hff6f;
  assign _zz_64 = 16'hff65;
  assign _zz__zz_A_15 = 16'h0001;
  assign _zz__zz_A_15_1 = 16'h0001;
  assign _zz__zz_A_15_2 = 16'h0001;
  assign _zz__zz_A_15_3 = 16'h0001;
  assign _zz__zz_A_15_4 = 16'h0001;
  assign _zz__zz_A_15_5 = 16'h0001;
  assign _zz__zz_A_15_6 = 16'h0001;
  assign _zz__zz_A_15_7 = 16'h0001;
  assign _zz__zz_A_15_8 = 16'h0001;
  assign _zz__zz_A_15_9 = 16'h0001;
  assign _zz__zz_A_15_10 = 16'h0001;
  assign _zz__zz_A_15_11 = 16'h0001;
  assign _zz__zz_A_15_12 = 16'h0001;
  assign _zz__zz_A_15_13 = 16'h0001;
  assign _zz__zz_A_15_14 = 16'h0001;
  assign _zz__zz_A_15_15 = 16'h0001;
  assign _zz__zz_A_15_16 = 16'h0001;
  assign _zz__zz_A_15_17 = 16'h0001;
  assign _zz__zz_A_15_18 = 16'h0001;
  assign _zz__zz_A_15_19 = 16'h0001;
  assign _zz__zz_A_15_20 = 16'h0001;
  assign _zz__zz_A_15_21 = 16'h0001;
  assign _zz__zz_A_15_22 = 16'h0001;
  assign _zz__zz_A_15_23 = 16'h0001;
  assign _zz__zz_A_15_24 = 16'h0001;
  assign _zz__zz_A_15_25 = 16'h0001;
  assign _zz__zz_A_15_26 = 16'h0001;
  assign _zz__zz_A_15_27 = 16'h0001;
  assign _zz__zz_A_15_28 = 16'h0001;
  assign _zz__zz_A_15_29 = 16'h0001;
  assign _zz__zz_A_15_30 = 16'h0001;
  assign _zz__zz_A_15_31 = 16'h0001;
  assign _zz__zz_dataOut_3 = _zz_dataOut_3_1;
  assign _zz_when_LeakyRelu_l157_3 = 16'h00ff;
  assign _zz__zz_A_17 = (_zz_when_LeakyRelu_l101_8 >>> 17);
  assign _zz__zz_A_17_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_4_1 = 4'b0000;
  assign _zz_65 = 16'hfffb;
  assign _zz_66 = 16'hfff1;
  assign _zz_67 = 16'hffe7;
  assign _zz_68 = 16'hffdd;
  assign _zz_69 = 16'hffd3;
  assign _zz_70 = 16'hffc9;
  assign _zz_71 = 16'hffbf;
  assign _zz_72 = 16'hffb5;
  assign _zz_73 = 16'hffab;
  assign _zz_74 = 16'hffa1;
  assign _zz_75 = 16'hff97;
  assign _zz_76 = 16'hff8d;
  assign _zz_77 = 16'hff83;
  assign _zz_78 = 16'hff79;
  assign _zz_79 = 16'hff6f;
  assign _zz_80 = 16'hff65;
  assign _zz__zz_A_19 = 16'h0001;
  assign _zz__zz_A_19_1 = 16'h0001;
  assign _zz__zz_A_19_2 = 16'h0001;
  assign _zz__zz_A_19_3 = 16'h0001;
  assign _zz__zz_A_19_4 = 16'h0001;
  assign _zz__zz_A_19_5 = 16'h0001;
  assign _zz__zz_A_19_6 = 16'h0001;
  assign _zz__zz_A_19_7 = 16'h0001;
  assign _zz__zz_A_19_8 = 16'h0001;
  assign _zz__zz_A_19_9 = 16'h0001;
  assign _zz__zz_A_19_10 = 16'h0001;
  assign _zz__zz_A_19_11 = 16'h0001;
  assign _zz__zz_A_19_12 = 16'h0001;
  assign _zz__zz_A_19_13 = 16'h0001;
  assign _zz__zz_A_19_14 = 16'h0001;
  assign _zz__zz_A_19_15 = 16'h0001;
  assign _zz__zz_A_19_16 = 16'h0001;
  assign _zz__zz_A_19_17 = 16'h0001;
  assign _zz__zz_A_19_18 = 16'h0001;
  assign _zz__zz_A_19_19 = 16'h0001;
  assign _zz__zz_A_19_20 = 16'h0001;
  assign _zz__zz_A_19_21 = 16'h0001;
  assign _zz__zz_A_19_22 = 16'h0001;
  assign _zz__zz_A_19_23 = 16'h0001;
  assign _zz__zz_A_19_24 = 16'h0001;
  assign _zz__zz_A_19_25 = 16'h0001;
  assign _zz__zz_A_19_26 = 16'h0001;
  assign _zz__zz_A_19_27 = 16'h0001;
  assign _zz__zz_A_19_28 = 16'h0001;
  assign _zz__zz_A_19_29 = 16'h0001;
  assign _zz__zz_A_19_30 = 16'h0001;
  assign _zz__zz_A_19_31 = 16'h0001;
  assign _zz__zz_dataOut_4 = _zz_dataOut_4_1;
  assign _zz_when_LeakyRelu_l157_4 = 16'h00ff;
  assign _zz__zz_A_21 = (_zz_when_LeakyRelu_l101_10 >>> 17);
  assign _zz__zz_A_21_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_5_1 = 4'b0000;
  assign _zz_81 = 16'hfffb;
  assign _zz_82 = 16'hfff1;
  assign _zz_83 = 16'hffe7;
  assign _zz_84 = 16'hffdd;
  assign _zz_85 = 16'hffd3;
  assign _zz_86 = 16'hffc9;
  assign _zz_87 = 16'hffbf;
  assign _zz_88 = 16'hffb5;
  assign _zz_89 = 16'hffab;
  assign _zz_90 = 16'hffa1;
  assign _zz_91 = 16'hff97;
  assign _zz_92 = 16'hff8d;
  assign _zz_93 = 16'hff83;
  assign _zz_94 = 16'hff79;
  assign _zz_95 = 16'hff6f;
  assign _zz_96 = 16'hff65;
  assign _zz__zz_A_23 = 16'h0001;
  assign _zz__zz_A_23_1 = 16'h0001;
  assign _zz__zz_A_23_2 = 16'h0001;
  assign _zz__zz_A_23_3 = 16'h0001;
  assign _zz__zz_A_23_4 = 16'h0001;
  assign _zz__zz_A_23_5 = 16'h0001;
  assign _zz__zz_A_23_6 = 16'h0001;
  assign _zz__zz_A_23_7 = 16'h0001;
  assign _zz__zz_A_23_8 = 16'h0001;
  assign _zz__zz_A_23_9 = 16'h0001;
  assign _zz__zz_A_23_10 = 16'h0001;
  assign _zz__zz_A_23_11 = 16'h0001;
  assign _zz__zz_A_23_12 = 16'h0001;
  assign _zz__zz_A_23_13 = 16'h0001;
  assign _zz__zz_A_23_14 = 16'h0001;
  assign _zz__zz_A_23_15 = 16'h0001;
  assign _zz__zz_A_23_16 = 16'h0001;
  assign _zz__zz_A_23_17 = 16'h0001;
  assign _zz__zz_A_23_18 = 16'h0001;
  assign _zz__zz_A_23_19 = 16'h0001;
  assign _zz__zz_A_23_20 = 16'h0001;
  assign _zz__zz_A_23_21 = 16'h0001;
  assign _zz__zz_A_23_22 = 16'h0001;
  assign _zz__zz_A_23_23 = 16'h0001;
  assign _zz__zz_A_23_24 = 16'h0001;
  assign _zz__zz_A_23_25 = 16'h0001;
  assign _zz__zz_A_23_26 = 16'h0001;
  assign _zz__zz_A_23_27 = 16'h0001;
  assign _zz__zz_A_23_28 = 16'h0001;
  assign _zz__zz_A_23_29 = 16'h0001;
  assign _zz__zz_A_23_30 = 16'h0001;
  assign _zz__zz_A_23_31 = 16'h0001;
  assign _zz__zz_dataOut_5 = _zz_dataOut_5_1;
  assign _zz_when_LeakyRelu_l157_5 = 16'h00ff;
  assign _zz__zz_A_25 = (_zz_when_LeakyRelu_l101_12 >>> 17);
  assign _zz__zz_A_25_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_6_1 = 4'b0000;
  assign _zz_97 = 16'hfffb;
  assign _zz_98 = 16'hfff1;
  assign _zz_99 = 16'hffe7;
  assign _zz_100 = 16'hffdd;
  assign _zz_101 = 16'hffd3;
  assign _zz_102 = 16'hffc9;
  assign _zz_103 = 16'hffbf;
  assign _zz_104 = 16'hffb5;
  assign _zz_105 = 16'hffab;
  assign _zz_106 = 16'hffa1;
  assign _zz_107 = 16'hff97;
  assign _zz_108 = 16'hff8d;
  assign _zz_109 = 16'hff83;
  assign _zz_110 = 16'hff79;
  assign _zz_111 = 16'hff6f;
  assign _zz_112 = 16'hff65;
  assign _zz__zz_A_27 = 16'h0001;
  assign _zz__zz_A_27_1 = 16'h0001;
  assign _zz__zz_A_27_2 = 16'h0001;
  assign _zz__zz_A_27_3 = 16'h0001;
  assign _zz__zz_A_27_4 = 16'h0001;
  assign _zz__zz_A_27_5 = 16'h0001;
  assign _zz__zz_A_27_6 = 16'h0001;
  assign _zz__zz_A_27_7 = 16'h0001;
  assign _zz__zz_A_27_8 = 16'h0001;
  assign _zz__zz_A_27_9 = 16'h0001;
  assign _zz__zz_A_27_10 = 16'h0001;
  assign _zz__zz_A_27_11 = 16'h0001;
  assign _zz__zz_A_27_12 = 16'h0001;
  assign _zz__zz_A_27_13 = 16'h0001;
  assign _zz__zz_A_27_14 = 16'h0001;
  assign _zz__zz_A_27_15 = 16'h0001;
  assign _zz__zz_A_27_16 = 16'h0001;
  assign _zz__zz_A_27_17 = 16'h0001;
  assign _zz__zz_A_27_18 = 16'h0001;
  assign _zz__zz_A_27_19 = 16'h0001;
  assign _zz__zz_A_27_20 = 16'h0001;
  assign _zz__zz_A_27_21 = 16'h0001;
  assign _zz__zz_A_27_22 = 16'h0001;
  assign _zz__zz_A_27_23 = 16'h0001;
  assign _zz__zz_A_27_24 = 16'h0001;
  assign _zz__zz_A_27_25 = 16'h0001;
  assign _zz__zz_A_27_26 = 16'h0001;
  assign _zz__zz_A_27_27 = 16'h0001;
  assign _zz__zz_A_27_28 = 16'h0001;
  assign _zz__zz_A_27_29 = 16'h0001;
  assign _zz__zz_A_27_30 = 16'h0001;
  assign _zz__zz_A_27_31 = 16'h0001;
  assign _zz__zz_dataOut_6 = _zz_dataOut_6_1;
  assign _zz_when_LeakyRelu_l157_6 = 16'h00ff;
  assign _zz__zz_A_29 = (_zz_when_LeakyRelu_l101_14 >>> 17);
  assign _zz__zz_A_29_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_7_1 = 4'b0000;
  assign _zz_113 = 16'hfffb;
  assign _zz_114 = 16'hfff1;
  assign _zz_115 = 16'hffe7;
  assign _zz_116 = 16'hffdd;
  assign _zz_117 = 16'hffd3;
  assign _zz_118 = 16'hffc9;
  assign _zz_119 = 16'hffbf;
  assign _zz_120 = 16'hffb5;
  assign _zz_121 = 16'hffab;
  assign _zz_122 = 16'hffa1;
  assign _zz_123 = 16'hff97;
  assign _zz_124 = 16'hff8d;
  assign _zz_125 = 16'hff83;
  assign _zz_126 = 16'hff79;
  assign _zz_127 = 16'hff6f;
  assign _zz_128 = 16'hff65;
  assign _zz__zz_A_31 = 16'h0001;
  assign _zz__zz_A_31_1 = 16'h0001;
  assign _zz__zz_A_31_2 = 16'h0001;
  assign _zz__zz_A_31_3 = 16'h0001;
  assign _zz__zz_A_31_4 = 16'h0001;
  assign _zz__zz_A_31_5 = 16'h0001;
  assign _zz__zz_A_31_6 = 16'h0001;
  assign _zz__zz_A_31_7 = 16'h0001;
  assign _zz__zz_A_31_8 = 16'h0001;
  assign _zz__zz_A_31_9 = 16'h0001;
  assign _zz__zz_A_31_10 = 16'h0001;
  assign _zz__zz_A_31_11 = 16'h0001;
  assign _zz__zz_A_31_12 = 16'h0001;
  assign _zz__zz_A_31_13 = 16'h0001;
  assign _zz__zz_A_31_14 = 16'h0001;
  assign _zz__zz_A_31_15 = 16'h0001;
  assign _zz__zz_A_31_16 = 16'h0001;
  assign _zz__zz_A_31_17 = 16'h0001;
  assign _zz__zz_A_31_18 = 16'h0001;
  assign _zz__zz_A_31_19 = 16'h0001;
  assign _zz__zz_A_31_20 = 16'h0001;
  assign _zz__zz_A_31_21 = 16'h0001;
  assign _zz__zz_A_31_22 = 16'h0001;
  assign _zz__zz_A_31_23 = 16'h0001;
  assign _zz__zz_A_31_24 = 16'h0001;
  assign _zz__zz_A_31_25 = 16'h0001;
  assign _zz__zz_A_31_26 = 16'h0001;
  assign _zz__zz_A_31_27 = 16'h0001;
  assign _zz__zz_A_31_28 = 16'h0001;
  assign _zz__zz_A_31_29 = 16'h0001;
  assign _zz__zz_A_31_30 = 16'h0001;
  assign _zz__zz_A_31_31 = 16'h0001;
  assign _zz__zz_dataOut_7 = _zz_dataOut_7_1;
  assign _zz_when_LeakyRelu_l157_7 = 16'h00ff;
  assign _zz__zz_A_33 = (_zz_when_LeakyRelu_l101_16 >>> 17);
  assign _zz__zz_A_33_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_8_1 = 4'b0000;
  assign _zz_129 = 16'hfffb;
  assign _zz_130 = 16'hfff1;
  assign _zz_131 = 16'hffe7;
  assign _zz_132 = 16'hffdd;
  assign _zz_133 = 16'hffd3;
  assign _zz_134 = 16'hffc9;
  assign _zz_135 = 16'hffbf;
  assign _zz_136 = 16'hffb5;
  assign _zz_137 = 16'hffab;
  assign _zz_138 = 16'hffa1;
  assign _zz_139 = 16'hff97;
  assign _zz_140 = 16'hff8d;
  assign _zz_141 = 16'hff83;
  assign _zz_142 = 16'hff79;
  assign _zz_143 = 16'hff6f;
  assign _zz_144 = 16'hff65;
  assign _zz__zz_A_35 = 16'h0001;
  assign _zz__zz_A_35_1 = 16'h0001;
  assign _zz__zz_A_35_2 = 16'h0001;
  assign _zz__zz_A_35_3 = 16'h0001;
  assign _zz__zz_A_35_4 = 16'h0001;
  assign _zz__zz_A_35_5 = 16'h0001;
  assign _zz__zz_A_35_6 = 16'h0001;
  assign _zz__zz_A_35_7 = 16'h0001;
  assign _zz__zz_A_35_8 = 16'h0001;
  assign _zz__zz_A_35_9 = 16'h0001;
  assign _zz__zz_A_35_10 = 16'h0001;
  assign _zz__zz_A_35_11 = 16'h0001;
  assign _zz__zz_A_35_12 = 16'h0001;
  assign _zz__zz_A_35_13 = 16'h0001;
  assign _zz__zz_A_35_14 = 16'h0001;
  assign _zz__zz_A_35_15 = 16'h0001;
  assign _zz__zz_A_35_16 = 16'h0001;
  assign _zz__zz_A_35_17 = 16'h0001;
  assign _zz__zz_A_35_18 = 16'h0001;
  assign _zz__zz_A_35_19 = 16'h0001;
  assign _zz__zz_A_35_20 = 16'h0001;
  assign _zz__zz_A_35_21 = 16'h0001;
  assign _zz__zz_A_35_22 = 16'h0001;
  assign _zz__zz_A_35_23 = 16'h0001;
  assign _zz__zz_A_35_24 = 16'h0001;
  assign _zz__zz_A_35_25 = 16'h0001;
  assign _zz__zz_A_35_26 = 16'h0001;
  assign _zz__zz_A_35_27 = 16'h0001;
  assign _zz__zz_A_35_28 = 16'h0001;
  assign _zz__zz_A_35_29 = 16'h0001;
  assign _zz__zz_A_35_30 = 16'h0001;
  assign _zz__zz_A_35_31 = 16'h0001;
  assign _zz__zz_dataOut_8 = _zz_dataOut_8_1;
  assign _zz_when_LeakyRelu_l157_8 = 16'h00ff;
  assign _zz__zz_A_37 = (_zz_when_LeakyRelu_l101_18 >>> 17);
  assign _zz__zz_A_37_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_9_1 = 4'b0000;
  assign _zz_145 = 16'hfffb;
  assign _zz_146 = 16'hfff1;
  assign _zz_147 = 16'hffe7;
  assign _zz_148 = 16'hffdd;
  assign _zz_149 = 16'hffd3;
  assign _zz_150 = 16'hffc9;
  assign _zz_151 = 16'hffbf;
  assign _zz_152 = 16'hffb5;
  assign _zz_153 = 16'hffab;
  assign _zz_154 = 16'hffa1;
  assign _zz_155 = 16'hff97;
  assign _zz_156 = 16'hff8d;
  assign _zz_157 = 16'hff83;
  assign _zz_158 = 16'hff79;
  assign _zz_159 = 16'hff6f;
  assign _zz_160 = 16'hff65;
  assign _zz__zz_A_39 = 16'h0001;
  assign _zz__zz_A_39_1 = 16'h0001;
  assign _zz__zz_A_39_2 = 16'h0001;
  assign _zz__zz_A_39_3 = 16'h0001;
  assign _zz__zz_A_39_4 = 16'h0001;
  assign _zz__zz_A_39_5 = 16'h0001;
  assign _zz__zz_A_39_6 = 16'h0001;
  assign _zz__zz_A_39_7 = 16'h0001;
  assign _zz__zz_A_39_8 = 16'h0001;
  assign _zz__zz_A_39_9 = 16'h0001;
  assign _zz__zz_A_39_10 = 16'h0001;
  assign _zz__zz_A_39_11 = 16'h0001;
  assign _zz__zz_A_39_12 = 16'h0001;
  assign _zz__zz_A_39_13 = 16'h0001;
  assign _zz__zz_A_39_14 = 16'h0001;
  assign _zz__zz_A_39_15 = 16'h0001;
  assign _zz__zz_A_39_16 = 16'h0001;
  assign _zz__zz_A_39_17 = 16'h0001;
  assign _zz__zz_A_39_18 = 16'h0001;
  assign _zz__zz_A_39_19 = 16'h0001;
  assign _zz__zz_A_39_20 = 16'h0001;
  assign _zz__zz_A_39_21 = 16'h0001;
  assign _zz__zz_A_39_22 = 16'h0001;
  assign _zz__zz_A_39_23 = 16'h0001;
  assign _zz__zz_A_39_24 = 16'h0001;
  assign _zz__zz_A_39_25 = 16'h0001;
  assign _zz__zz_A_39_26 = 16'h0001;
  assign _zz__zz_A_39_27 = 16'h0001;
  assign _zz__zz_A_39_28 = 16'h0001;
  assign _zz__zz_A_39_29 = 16'h0001;
  assign _zz__zz_A_39_30 = 16'h0001;
  assign _zz__zz_A_39_31 = 16'h0001;
  assign _zz__zz_dataOut_9 = _zz_dataOut_9_1;
  assign _zz_when_LeakyRelu_l157_9 = 16'h00ff;
  assign _zz__zz_A_41 = (_zz_when_LeakyRelu_l101_20 >>> 17);
  assign _zz__zz_A_41_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_10_1 = 4'b0000;
  assign _zz_161 = 16'hfffb;
  assign _zz_162 = 16'hfff1;
  assign _zz_163 = 16'hffe7;
  assign _zz_164 = 16'hffdd;
  assign _zz_165 = 16'hffd3;
  assign _zz_166 = 16'hffc9;
  assign _zz_167 = 16'hffbf;
  assign _zz_168 = 16'hffb5;
  assign _zz_169 = 16'hffab;
  assign _zz_170 = 16'hffa1;
  assign _zz_171 = 16'hff97;
  assign _zz_172 = 16'hff8d;
  assign _zz_173 = 16'hff83;
  assign _zz_174 = 16'hff79;
  assign _zz_175 = 16'hff6f;
  assign _zz_176 = 16'hff65;
  assign _zz__zz_A_43 = 16'h0001;
  assign _zz__zz_A_43_1 = 16'h0001;
  assign _zz__zz_A_43_2 = 16'h0001;
  assign _zz__zz_A_43_3 = 16'h0001;
  assign _zz__zz_A_43_4 = 16'h0001;
  assign _zz__zz_A_43_5 = 16'h0001;
  assign _zz__zz_A_43_6 = 16'h0001;
  assign _zz__zz_A_43_7 = 16'h0001;
  assign _zz__zz_A_43_8 = 16'h0001;
  assign _zz__zz_A_43_9 = 16'h0001;
  assign _zz__zz_A_43_10 = 16'h0001;
  assign _zz__zz_A_43_11 = 16'h0001;
  assign _zz__zz_A_43_12 = 16'h0001;
  assign _zz__zz_A_43_13 = 16'h0001;
  assign _zz__zz_A_43_14 = 16'h0001;
  assign _zz__zz_A_43_15 = 16'h0001;
  assign _zz__zz_A_43_16 = 16'h0001;
  assign _zz__zz_A_43_17 = 16'h0001;
  assign _zz__zz_A_43_18 = 16'h0001;
  assign _zz__zz_A_43_19 = 16'h0001;
  assign _zz__zz_A_43_20 = 16'h0001;
  assign _zz__zz_A_43_21 = 16'h0001;
  assign _zz__zz_A_43_22 = 16'h0001;
  assign _zz__zz_A_43_23 = 16'h0001;
  assign _zz__zz_A_43_24 = 16'h0001;
  assign _zz__zz_A_43_25 = 16'h0001;
  assign _zz__zz_A_43_26 = 16'h0001;
  assign _zz__zz_A_43_27 = 16'h0001;
  assign _zz__zz_A_43_28 = 16'h0001;
  assign _zz__zz_A_43_29 = 16'h0001;
  assign _zz__zz_A_43_30 = 16'h0001;
  assign _zz__zz_A_43_31 = 16'h0001;
  assign _zz__zz_dataOut_10 = _zz_dataOut_10_1;
  assign _zz_when_LeakyRelu_l157_10 = 16'h00ff;
  assign _zz__zz_A_45 = (_zz_when_LeakyRelu_l101_22 >>> 17);
  assign _zz__zz_A_45_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_11_1 = 4'b0000;
  assign _zz_177 = 16'hfffb;
  assign _zz_178 = 16'hfff1;
  assign _zz_179 = 16'hffe7;
  assign _zz_180 = 16'hffdd;
  assign _zz_181 = 16'hffd3;
  assign _zz_182 = 16'hffc9;
  assign _zz_183 = 16'hffbf;
  assign _zz_184 = 16'hffb5;
  assign _zz_185 = 16'hffab;
  assign _zz_186 = 16'hffa1;
  assign _zz_187 = 16'hff97;
  assign _zz_188 = 16'hff8d;
  assign _zz_189 = 16'hff83;
  assign _zz_190 = 16'hff79;
  assign _zz_191 = 16'hff6f;
  assign _zz_192 = 16'hff65;
  assign _zz__zz_A_47 = 16'h0001;
  assign _zz__zz_A_47_1 = 16'h0001;
  assign _zz__zz_A_47_2 = 16'h0001;
  assign _zz__zz_A_47_3 = 16'h0001;
  assign _zz__zz_A_47_4 = 16'h0001;
  assign _zz__zz_A_47_5 = 16'h0001;
  assign _zz__zz_A_47_6 = 16'h0001;
  assign _zz__zz_A_47_7 = 16'h0001;
  assign _zz__zz_A_47_8 = 16'h0001;
  assign _zz__zz_A_47_9 = 16'h0001;
  assign _zz__zz_A_47_10 = 16'h0001;
  assign _zz__zz_A_47_11 = 16'h0001;
  assign _zz__zz_A_47_12 = 16'h0001;
  assign _zz__zz_A_47_13 = 16'h0001;
  assign _zz__zz_A_47_14 = 16'h0001;
  assign _zz__zz_A_47_15 = 16'h0001;
  assign _zz__zz_A_47_16 = 16'h0001;
  assign _zz__zz_A_47_17 = 16'h0001;
  assign _zz__zz_A_47_18 = 16'h0001;
  assign _zz__zz_A_47_19 = 16'h0001;
  assign _zz__zz_A_47_20 = 16'h0001;
  assign _zz__zz_A_47_21 = 16'h0001;
  assign _zz__zz_A_47_22 = 16'h0001;
  assign _zz__zz_A_47_23 = 16'h0001;
  assign _zz__zz_A_47_24 = 16'h0001;
  assign _zz__zz_A_47_25 = 16'h0001;
  assign _zz__zz_A_47_26 = 16'h0001;
  assign _zz__zz_A_47_27 = 16'h0001;
  assign _zz__zz_A_47_28 = 16'h0001;
  assign _zz__zz_A_47_29 = 16'h0001;
  assign _zz__zz_A_47_30 = 16'h0001;
  assign _zz__zz_A_47_31 = 16'h0001;
  assign _zz__zz_dataOut_11 = _zz_dataOut_11_1;
  assign _zz_when_LeakyRelu_l157_11 = 16'h00ff;
  assign _zz__zz_A_49 = (_zz_when_LeakyRelu_l101_24 >>> 17);
  assign _zz__zz_A_49_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_12_1 = 4'b0000;
  assign _zz_193 = 16'hfffb;
  assign _zz_194 = 16'hfff1;
  assign _zz_195 = 16'hffe7;
  assign _zz_196 = 16'hffdd;
  assign _zz_197 = 16'hffd3;
  assign _zz_198 = 16'hffc9;
  assign _zz_199 = 16'hffbf;
  assign _zz_200 = 16'hffb5;
  assign _zz_201 = 16'hffab;
  assign _zz_202 = 16'hffa1;
  assign _zz_203 = 16'hff97;
  assign _zz_204 = 16'hff8d;
  assign _zz_205 = 16'hff83;
  assign _zz_206 = 16'hff79;
  assign _zz_207 = 16'hff6f;
  assign _zz_208 = 16'hff65;
  assign _zz__zz_A_51 = 16'h0001;
  assign _zz__zz_A_51_1 = 16'h0001;
  assign _zz__zz_A_51_2 = 16'h0001;
  assign _zz__zz_A_51_3 = 16'h0001;
  assign _zz__zz_A_51_4 = 16'h0001;
  assign _zz__zz_A_51_5 = 16'h0001;
  assign _zz__zz_A_51_6 = 16'h0001;
  assign _zz__zz_A_51_7 = 16'h0001;
  assign _zz__zz_A_51_8 = 16'h0001;
  assign _zz__zz_A_51_9 = 16'h0001;
  assign _zz__zz_A_51_10 = 16'h0001;
  assign _zz__zz_A_51_11 = 16'h0001;
  assign _zz__zz_A_51_12 = 16'h0001;
  assign _zz__zz_A_51_13 = 16'h0001;
  assign _zz__zz_A_51_14 = 16'h0001;
  assign _zz__zz_A_51_15 = 16'h0001;
  assign _zz__zz_A_51_16 = 16'h0001;
  assign _zz__zz_A_51_17 = 16'h0001;
  assign _zz__zz_A_51_18 = 16'h0001;
  assign _zz__zz_A_51_19 = 16'h0001;
  assign _zz__zz_A_51_20 = 16'h0001;
  assign _zz__zz_A_51_21 = 16'h0001;
  assign _zz__zz_A_51_22 = 16'h0001;
  assign _zz__zz_A_51_23 = 16'h0001;
  assign _zz__zz_A_51_24 = 16'h0001;
  assign _zz__zz_A_51_25 = 16'h0001;
  assign _zz__zz_A_51_26 = 16'h0001;
  assign _zz__zz_A_51_27 = 16'h0001;
  assign _zz__zz_A_51_28 = 16'h0001;
  assign _zz__zz_A_51_29 = 16'h0001;
  assign _zz__zz_A_51_30 = 16'h0001;
  assign _zz__zz_A_51_31 = 16'h0001;
  assign _zz__zz_dataOut_12 = _zz_dataOut_12_1;
  assign _zz_when_LeakyRelu_l157_12 = 16'h00ff;
  assign _zz__zz_A_53 = (_zz_when_LeakyRelu_l101_26 >>> 17);
  assign _zz__zz_A_53_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_13_1 = 4'b0000;
  assign _zz_209 = 16'hfffb;
  assign _zz_210 = 16'hfff1;
  assign _zz_211 = 16'hffe7;
  assign _zz_212 = 16'hffdd;
  assign _zz_213 = 16'hffd3;
  assign _zz_214 = 16'hffc9;
  assign _zz_215 = 16'hffbf;
  assign _zz_216 = 16'hffb5;
  assign _zz_217 = 16'hffab;
  assign _zz_218 = 16'hffa1;
  assign _zz_219 = 16'hff97;
  assign _zz_220 = 16'hff8d;
  assign _zz_221 = 16'hff83;
  assign _zz_222 = 16'hff79;
  assign _zz_223 = 16'hff6f;
  assign _zz_224 = 16'hff65;
  assign _zz__zz_A_55 = 16'h0001;
  assign _zz__zz_A_55_1 = 16'h0001;
  assign _zz__zz_A_55_2 = 16'h0001;
  assign _zz__zz_A_55_3 = 16'h0001;
  assign _zz__zz_A_55_4 = 16'h0001;
  assign _zz__zz_A_55_5 = 16'h0001;
  assign _zz__zz_A_55_6 = 16'h0001;
  assign _zz__zz_A_55_7 = 16'h0001;
  assign _zz__zz_A_55_8 = 16'h0001;
  assign _zz__zz_A_55_9 = 16'h0001;
  assign _zz__zz_A_55_10 = 16'h0001;
  assign _zz__zz_A_55_11 = 16'h0001;
  assign _zz__zz_A_55_12 = 16'h0001;
  assign _zz__zz_A_55_13 = 16'h0001;
  assign _zz__zz_A_55_14 = 16'h0001;
  assign _zz__zz_A_55_15 = 16'h0001;
  assign _zz__zz_A_55_16 = 16'h0001;
  assign _zz__zz_A_55_17 = 16'h0001;
  assign _zz__zz_A_55_18 = 16'h0001;
  assign _zz__zz_A_55_19 = 16'h0001;
  assign _zz__zz_A_55_20 = 16'h0001;
  assign _zz__zz_A_55_21 = 16'h0001;
  assign _zz__zz_A_55_22 = 16'h0001;
  assign _zz__zz_A_55_23 = 16'h0001;
  assign _zz__zz_A_55_24 = 16'h0001;
  assign _zz__zz_A_55_25 = 16'h0001;
  assign _zz__zz_A_55_26 = 16'h0001;
  assign _zz__zz_A_55_27 = 16'h0001;
  assign _zz__zz_A_55_28 = 16'h0001;
  assign _zz__zz_A_55_29 = 16'h0001;
  assign _zz__zz_A_55_30 = 16'h0001;
  assign _zz__zz_A_55_31 = 16'h0001;
  assign _zz__zz_dataOut_13 = _zz_dataOut_13_1;
  assign _zz_when_LeakyRelu_l157_13 = 16'h00ff;
  assign _zz__zz_A_57 = (_zz_when_LeakyRelu_l101_28 >>> 17);
  assign _zz__zz_A_57_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_14_1 = 4'b0000;
  assign _zz_225 = 16'hfffb;
  assign _zz_226 = 16'hfff1;
  assign _zz_227 = 16'hffe7;
  assign _zz_228 = 16'hffdd;
  assign _zz_229 = 16'hffd3;
  assign _zz_230 = 16'hffc9;
  assign _zz_231 = 16'hffbf;
  assign _zz_232 = 16'hffb5;
  assign _zz_233 = 16'hffab;
  assign _zz_234 = 16'hffa1;
  assign _zz_235 = 16'hff97;
  assign _zz_236 = 16'hff8d;
  assign _zz_237 = 16'hff83;
  assign _zz_238 = 16'hff79;
  assign _zz_239 = 16'hff6f;
  assign _zz_240 = 16'hff65;
  assign _zz__zz_A_59 = 16'h0001;
  assign _zz__zz_A_59_1 = 16'h0001;
  assign _zz__zz_A_59_2 = 16'h0001;
  assign _zz__zz_A_59_3 = 16'h0001;
  assign _zz__zz_A_59_4 = 16'h0001;
  assign _zz__zz_A_59_5 = 16'h0001;
  assign _zz__zz_A_59_6 = 16'h0001;
  assign _zz__zz_A_59_7 = 16'h0001;
  assign _zz__zz_A_59_8 = 16'h0001;
  assign _zz__zz_A_59_9 = 16'h0001;
  assign _zz__zz_A_59_10 = 16'h0001;
  assign _zz__zz_A_59_11 = 16'h0001;
  assign _zz__zz_A_59_12 = 16'h0001;
  assign _zz__zz_A_59_13 = 16'h0001;
  assign _zz__zz_A_59_14 = 16'h0001;
  assign _zz__zz_A_59_15 = 16'h0001;
  assign _zz__zz_A_59_16 = 16'h0001;
  assign _zz__zz_A_59_17 = 16'h0001;
  assign _zz__zz_A_59_18 = 16'h0001;
  assign _zz__zz_A_59_19 = 16'h0001;
  assign _zz__zz_A_59_20 = 16'h0001;
  assign _zz__zz_A_59_21 = 16'h0001;
  assign _zz__zz_A_59_22 = 16'h0001;
  assign _zz__zz_A_59_23 = 16'h0001;
  assign _zz__zz_A_59_24 = 16'h0001;
  assign _zz__zz_A_59_25 = 16'h0001;
  assign _zz__zz_A_59_26 = 16'h0001;
  assign _zz__zz_A_59_27 = 16'h0001;
  assign _zz__zz_A_59_28 = 16'h0001;
  assign _zz__zz_A_59_29 = 16'h0001;
  assign _zz__zz_A_59_30 = 16'h0001;
  assign _zz__zz_A_59_31 = 16'h0001;
  assign _zz__zz_dataOut_14 = _zz_dataOut_14_1;
  assign _zz_when_LeakyRelu_l157_14 = 16'h00ff;
  assign _zz__zz_A_61 = (_zz_when_LeakyRelu_l101_30 >>> 17);
  assign _zz__zz_A_61_1 = 15'h0001;
  assign _zz_when_LeakyRelu_l101_15_1 = 4'b0000;
  assign _zz_241 = 16'hfffb;
  assign _zz_242 = 16'hfff1;
  assign _zz_243 = 16'hffe7;
  assign _zz_244 = 16'hffdd;
  assign _zz_245 = 16'hffd3;
  assign _zz_246 = 16'hffc9;
  assign _zz_247 = 16'hffbf;
  assign _zz_248 = 16'hffb5;
  assign _zz_249 = 16'hffab;
  assign _zz_250 = 16'hffa1;
  assign _zz_251 = 16'hff97;
  assign _zz_252 = 16'hff8d;
  assign _zz_253 = 16'hff83;
  assign _zz_254 = 16'hff79;
  assign _zz_255 = 16'hff6f;
  assign _zz_256 = 16'hff65;
  assign _zz__zz_A_63 = 16'h0001;
  assign _zz__zz_A_63_1 = 16'h0001;
  assign _zz__zz_A_63_2 = 16'h0001;
  assign _zz__zz_A_63_3 = 16'h0001;
  assign _zz__zz_A_63_4 = 16'h0001;
  assign _zz__zz_A_63_5 = 16'h0001;
  assign _zz__zz_A_63_6 = 16'h0001;
  assign _zz__zz_A_63_7 = 16'h0001;
  assign _zz__zz_A_63_8 = 16'h0001;
  assign _zz__zz_A_63_9 = 16'h0001;
  assign _zz__zz_A_63_10 = 16'h0001;
  assign _zz__zz_A_63_11 = 16'h0001;
  assign _zz__zz_A_63_12 = 16'h0001;
  assign _zz__zz_A_63_13 = 16'h0001;
  assign _zz__zz_A_63_14 = 16'h0001;
  assign _zz__zz_A_63_15 = 16'h0001;
  assign _zz__zz_A_63_16 = 16'h0001;
  assign _zz__zz_A_63_17 = 16'h0001;
  assign _zz__zz_A_63_18 = 16'h0001;
  assign _zz__zz_A_63_19 = 16'h0001;
  assign _zz__zz_A_63_20 = 16'h0001;
  assign _zz__zz_A_63_21 = 16'h0001;
  assign _zz__zz_A_63_22 = 16'h0001;
  assign _zz__zz_A_63_23 = 16'h0001;
  assign _zz__zz_A_63_24 = 16'h0001;
  assign _zz__zz_A_63_25 = 16'h0001;
  assign _zz__zz_A_63_26 = 16'h0001;
  assign _zz__zz_A_63_27 = 16'h0001;
  assign _zz__zz_A_63_28 = 16'h0001;
  assign _zz__zz_A_63_29 = 16'h0001;
  assign _zz__zz_A_63_30 = 16'h0001;
  assign _zz__zz_A_63_31 = 16'h0001;
  assign _zz__zz_dataOut_15 = _zz_dataOut_15_1;
  assign _zz_when_LeakyRelu_l157_15 = 16'h00ff;
  leakySubZ3 addSub (
    .A   (addSub_A[15:0]), //i
    .B   (quanZero[7:0] ), //i
    .S   (addSub_S[15:0]), //o
    .CLK (clk           )  //i
  );
  leakyReluMul mul (
    .A   (_zz_when_LeakyRelu_l100[15:0]), //i
    .B   (leaky[15:0]                  ), //i
    .P   (mul_P[31:0]                  ), //o
    .CLK (clk                          )  //i
  );
  leakyAddZ3 addSub_1 (
    .A   (_zz_A_3[15:0]   ), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_1_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakySubZ3 addSub_2 (
    .A   (addSub_2_A[15:0]), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_2_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakyReluMul mul_1 (
    .A   (_zz_when_LeakyRelu_l100_4[15:0]), //i
    .B   (leaky[15:0]                    ), //i
    .P   (mul_1_P[31:0]                  ), //o
    .CLK (clk                            )  //i
  );
  leakyAddZ3 addSub_3 (
    .A   (_zz_A_7[15:0]   ), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_3_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakySubZ3 addSub_4 (
    .A   (addSub_4_A[15:0]), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_4_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakyReluMul mul_2 (
    .A   (_zz_when_LeakyRelu_l100_8[15:0]), //i
    .B   (leaky[15:0]                    ), //i
    .P   (mul_2_P[31:0]                  ), //o
    .CLK (clk                            )  //i
  );
  leakyAddZ3 addSub_5 (
    .A   (_zz_A_11[15:0]  ), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_5_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakySubZ3 addSub_6 (
    .A   (addSub_6_A[15:0]), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_6_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakyReluMul mul_3 (
    .A   (_zz_when_LeakyRelu_l100_12[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_3_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_7 (
    .A   (_zz_A_15[15:0]  ), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_7_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakySubZ3 addSub_8 (
    .A   (addSub_8_A[15:0]), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_8_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakyReluMul mul_4 (
    .A   (_zz_when_LeakyRelu_l100_16[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_4_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_9 (
    .A   (_zz_A_19[15:0]  ), //i
    .B   (quanZero[7:0]   ), //i
    .S   (addSub_9_S[15:0]), //o
    .CLK (clk             )  //i
  );
  leakySubZ3 addSub_10 (
    .A   (addSub_10_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_10_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_5 (
    .A   (_zz_when_LeakyRelu_l100_20[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_5_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_11 (
    .A   (_zz_A_23[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_11_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_12 (
    .A   (addSub_12_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_12_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_6 (
    .A   (_zz_when_LeakyRelu_l100_24[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_6_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_13 (
    .A   (_zz_A_27[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_13_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_14 (
    .A   (addSub_14_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_14_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_7 (
    .A   (_zz_when_LeakyRelu_l100_28[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_7_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_15 (
    .A   (_zz_A_31[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_15_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_16 (
    .A   (addSub_16_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_16_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_8 (
    .A   (_zz_when_LeakyRelu_l100_32[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_8_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_17 (
    .A   (_zz_A_35[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_17_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_18 (
    .A   (addSub_18_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_18_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_9 (
    .A   (_zz_when_LeakyRelu_l100_36[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_9_P[31:0]                   ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_19 (
    .A   (_zz_A_39[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_19_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_20 (
    .A   (addSub_20_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_20_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_10 (
    .A   (_zz_when_LeakyRelu_l100_40[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_10_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_21 (
    .A   (_zz_A_43[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_21_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_22 (
    .A   (addSub_22_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_22_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_11 (
    .A   (_zz_when_LeakyRelu_l100_44[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_11_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_23 (
    .A   (_zz_A_47[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_23_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_24 (
    .A   (addSub_24_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_24_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_12 (
    .A   (_zz_when_LeakyRelu_l100_48[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_12_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_25 (
    .A   (_zz_A_51[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_25_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_26 (
    .A   (addSub_26_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_26_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_13 (
    .A   (_zz_when_LeakyRelu_l100_52[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_13_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_27 (
    .A   (_zz_A_55[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_27_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_28 (
    .A   (addSub_28_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_28_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_14 (
    .A   (_zz_when_LeakyRelu_l100_56[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_14_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_29 (
    .A   (_zz_A_59[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_29_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakySubZ3 addSub_30 (
    .A   (addSub_30_A[15:0]), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_30_S[15:0]), //o
    .CLK (clk              )  //i
  );
  leakyReluMul mul_15 (
    .A   (_zz_when_LeakyRelu_l100_60[15:0]), //i
    .B   (leaky[15:0]                     ), //i
    .P   (mul_15_P[31:0]                  ), //o
    .CLK (clk                             )  //i
  );
  leakyAddZ3 addSub_31 (
    .A   (_zz_A_63[15:0]   ), //i
    .B   (quanZero[7:0]    ), //i
    .S   (addSub_31_S[15:0]), //o
    .CLK (clk              )  //i
  );
  assign leaky = 16'h3333;
  assign addSub_A = {8'h0,dataIn_0};
  assign _zz_when_LeakyRelu_l100 = addSub_S;
  assign _zz_when_LeakyRelu_l101_1 = _zz_when_LeakyRelu_l101[16 : 13];
  assign _zz_A_1 = ($signed(_zz__zz_A_1) + $signed(_zz__zz_A_1_1));
  assign _zz_A_2 = (_zz_when_LeakyRelu_l101 >>> 17);
  assign _zz_when_LeakyRelu_l101 = mul_P;
  assign when_LeakyRelu_l100 = _zz_when_LeakyRelu_l100_3[15];
  assign when_LeakyRelu_l101 = ($signed(_zz_when_LeakyRelu_l101_1) == $signed(_zz_when_LeakyRelu_l101_32));
  assign when_LeakyRelu_l104 = _zz_when_LeakyRelu_l101[16];
  assign when_LeakyRelu_l110 = (4'b1000 < _zz_when_LeakyRelu_l101_1);
  assign when_LeakyRelu_l103 = _zz_when_LeakyRelu_l101[17];
  assign when_LeakyRelu_l127 = _zz_when_LeakyRelu_l100_3_regNext[15];
  assign when_LeakyRelu_l131 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_1 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_1 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_2 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_2 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_3 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_3 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_4 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_4 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_5 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_5 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_6 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_6 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_7 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_7 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_8 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_8 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_9 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_9 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_10 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_10 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_11 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_11 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_12 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_12 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_13 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_13 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_14 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_14 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_15 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_15 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_0_1 = addSub_1_S;
  assign when_LeakyRelu_l155 = _zz_dataOut_0_1[15];
  assign when_LeakyRelu_l157 = ($signed(_zz_when_LeakyRelu_l157) < $signed(_zz_dataOut_0_1));
  assign dataOut_0 = _zz_dataOut_0;
  assign addSub_2_A = {8'h0,dataIn_1};
  assign _zz_when_LeakyRelu_l100_4 = addSub_2_S;
  assign _zz_when_LeakyRelu_l101_3 = _zz_when_LeakyRelu_l101_2[16 : 13];
  assign _zz_A_5 = ($signed(_zz__zz_A_5) + $signed(_zz__zz_A_5_1));
  assign _zz_A_6 = (_zz_when_LeakyRelu_l101_2 >>> 17);
  assign _zz_when_LeakyRelu_l101_2 = mul_1_P;
  assign when_LeakyRelu_l100_1 = _zz_when_LeakyRelu_l100_7[15];
  assign when_LeakyRelu_l101_1 = ($signed(_zz_when_LeakyRelu_l101_3) == $signed(_zz_when_LeakyRelu_l101_1_1));
  assign when_LeakyRelu_l104_1 = _zz_when_LeakyRelu_l101_2[16];
  assign when_LeakyRelu_l110_1 = (4'b1000 < _zz_when_LeakyRelu_l101_3);
  assign when_LeakyRelu_l103_1 = _zz_when_LeakyRelu_l101_2[17];
  assign when_LeakyRelu_l127_1 = _zz_when_LeakyRelu_l100_7_regNext[15];
  assign when_LeakyRelu_l131_16 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_16 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_17 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_17 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_18 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_18 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_19 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_19 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_20 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_20 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_21 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_21 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_22 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_22 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_23 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_23 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_24 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_24 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_25 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_25 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_26 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_26 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_27 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_27 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_28 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_28 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_29 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_29 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_30 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_30 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_31 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_31 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_1_1 = addSub_3_S;
  assign when_LeakyRelu_l155_1 = _zz_dataOut_1_1[15];
  assign when_LeakyRelu_l157_1 = ($signed(_zz_when_LeakyRelu_l157_1) < $signed(_zz_dataOut_1_1));
  assign dataOut_1 = _zz_dataOut_1;
  assign addSub_4_A = {8'h0,dataIn_2};
  assign _zz_when_LeakyRelu_l100_8 = addSub_4_S;
  assign _zz_when_LeakyRelu_l101_5 = _zz_when_LeakyRelu_l101_4[16 : 13];
  assign _zz_A_9 = ($signed(_zz__zz_A_9) + $signed(_zz__zz_A_9_1));
  assign _zz_A_10 = (_zz_when_LeakyRelu_l101_4 >>> 17);
  assign _zz_when_LeakyRelu_l101_4 = mul_2_P;
  assign when_LeakyRelu_l100_2 = _zz_when_LeakyRelu_l100_11[15];
  assign when_LeakyRelu_l101_2 = ($signed(_zz_when_LeakyRelu_l101_5) == $signed(_zz_when_LeakyRelu_l101_2_1));
  assign when_LeakyRelu_l104_2 = _zz_when_LeakyRelu_l101_4[16];
  assign when_LeakyRelu_l110_2 = (4'b1000 < _zz_when_LeakyRelu_l101_5);
  assign when_LeakyRelu_l103_2 = _zz_when_LeakyRelu_l101_4[17];
  assign when_LeakyRelu_l127_2 = _zz_when_LeakyRelu_l100_11_regNext[15];
  assign when_LeakyRelu_l131_32 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_32 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_33 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_33 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_34 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_34 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_35 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_35 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_36 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_36 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_37 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_37 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_38 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_38 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_39 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_39 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_40 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_40 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_41 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_41 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_42 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_42 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_43 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_43 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_44 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_44 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_45 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_45 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_46 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_46 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_47 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_47 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_2_1 = addSub_5_S;
  assign when_LeakyRelu_l155_2 = _zz_dataOut_2_1[15];
  assign when_LeakyRelu_l157_2 = ($signed(_zz_when_LeakyRelu_l157_2) < $signed(_zz_dataOut_2_1));
  assign dataOut_2 = _zz_dataOut_2;
  assign addSub_6_A = {8'h0,dataIn_3};
  assign _zz_when_LeakyRelu_l100_12 = addSub_6_S;
  assign _zz_when_LeakyRelu_l101_7 = _zz_when_LeakyRelu_l101_6[16 : 13];
  assign _zz_A_13 = ($signed(_zz__zz_A_13) + $signed(_zz__zz_A_13_1));
  assign _zz_A_14 = (_zz_when_LeakyRelu_l101_6 >>> 17);
  assign _zz_when_LeakyRelu_l101_6 = mul_3_P;
  assign when_LeakyRelu_l100_3 = _zz_when_LeakyRelu_l100_15[15];
  assign when_LeakyRelu_l101_3 = ($signed(_zz_when_LeakyRelu_l101_7) == $signed(_zz_when_LeakyRelu_l101_3_1));
  assign when_LeakyRelu_l104_3 = _zz_when_LeakyRelu_l101_6[16];
  assign when_LeakyRelu_l110_3 = (4'b1000 < _zz_when_LeakyRelu_l101_7);
  assign when_LeakyRelu_l103_3 = _zz_when_LeakyRelu_l101_6[17];
  assign when_LeakyRelu_l127_3 = _zz_when_LeakyRelu_l100_15_regNext[15];
  assign when_LeakyRelu_l131_48 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_48 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_49 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_49 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_50 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_50 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_51 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_51 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_52 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_52 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_53 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_53 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_54 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_54 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_55 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_55 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_56 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_56 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_57 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_57 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_58 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_58 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_59 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_59 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_60 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_60 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_61 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_61 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_62 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_62 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_63 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_63 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_3_1 = addSub_7_S;
  assign when_LeakyRelu_l155_3 = _zz_dataOut_3_1[15];
  assign when_LeakyRelu_l157_3 = ($signed(_zz_when_LeakyRelu_l157_3) < $signed(_zz_dataOut_3_1));
  assign dataOut_3 = _zz_dataOut_3;
  assign addSub_8_A = {8'h0,dataIn_4};
  assign _zz_when_LeakyRelu_l100_16 = addSub_8_S;
  assign _zz_when_LeakyRelu_l101_9 = _zz_when_LeakyRelu_l101_8[16 : 13];
  assign _zz_A_17 = ($signed(_zz__zz_A_17) + $signed(_zz__zz_A_17_1));
  assign _zz_A_18 = (_zz_when_LeakyRelu_l101_8 >>> 17);
  assign _zz_when_LeakyRelu_l101_8 = mul_4_P;
  assign when_LeakyRelu_l100_4 = _zz_when_LeakyRelu_l100_19[15];
  assign when_LeakyRelu_l101_4 = ($signed(_zz_when_LeakyRelu_l101_9) == $signed(_zz_when_LeakyRelu_l101_4_1));
  assign when_LeakyRelu_l104_4 = _zz_when_LeakyRelu_l101_8[16];
  assign when_LeakyRelu_l110_4 = (4'b1000 < _zz_when_LeakyRelu_l101_9);
  assign when_LeakyRelu_l103_4 = _zz_when_LeakyRelu_l101_8[17];
  assign when_LeakyRelu_l127_4 = _zz_when_LeakyRelu_l100_19_regNext[15];
  assign when_LeakyRelu_l131_64 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_64 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_65 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_65 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_66 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_66 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_67 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_67 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_68 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_68 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_69 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_69 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_70 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_70 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_71 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_71 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_72 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_72 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_73 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_73 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_74 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_74 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_75 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_75 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_76 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_76 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_77 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_77 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_78 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_78 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_79 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_79 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_4_1 = addSub_9_S;
  assign when_LeakyRelu_l155_4 = _zz_dataOut_4_1[15];
  assign when_LeakyRelu_l157_4 = ($signed(_zz_when_LeakyRelu_l157_4) < $signed(_zz_dataOut_4_1));
  assign dataOut_4 = _zz_dataOut_4;
  assign addSub_10_A = {8'h0,dataIn_5};
  assign _zz_when_LeakyRelu_l100_20 = addSub_10_S;
  assign _zz_when_LeakyRelu_l101_11 = _zz_when_LeakyRelu_l101_10[16 : 13];
  assign _zz_A_21 = ($signed(_zz__zz_A_21) + $signed(_zz__zz_A_21_1));
  assign _zz_A_22 = (_zz_when_LeakyRelu_l101_10 >>> 17);
  assign _zz_when_LeakyRelu_l101_10 = mul_5_P;
  assign when_LeakyRelu_l100_5 = _zz_when_LeakyRelu_l100_23[15];
  assign when_LeakyRelu_l101_5 = ($signed(_zz_when_LeakyRelu_l101_11) == $signed(_zz_when_LeakyRelu_l101_5_1));
  assign when_LeakyRelu_l104_5 = _zz_when_LeakyRelu_l101_10[16];
  assign when_LeakyRelu_l110_5 = (4'b1000 < _zz_when_LeakyRelu_l101_11);
  assign when_LeakyRelu_l103_5 = _zz_when_LeakyRelu_l101_10[17];
  assign when_LeakyRelu_l127_5 = _zz_when_LeakyRelu_l100_23_regNext[15];
  assign when_LeakyRelu_l131_80 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_80 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_81 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_81 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_82 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_82 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_83 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_83 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_84 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_84 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_85 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_85 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_86 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_86 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_87 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_87 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_88 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_88 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_89 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_89 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_90 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_90 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_91 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_91 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_92 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_92 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_93 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_93 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_94 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_94 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_95 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_95 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_5_1 = addSub_11_S;
  assign when_LeakyRelu_l155_5 = _zz_dataOut_5_1[15];
  assign when_LeakyRelu_l157_5 = ($signed(_zz_when_LeakyRelu_l157_5) < $signed(_zz_dataOut_5_1));
  assign dataOut_5 = _zz_dataOut_5;
  assign addSub_12_A = {8'h0,dataIn_6};
  assign _zz_when_LeakyRelu_l100_24 = addSub_12_S;
  assign _zz_when_LeakyRelu_l101_13 = _zz_when_LeakyRelu_l101_12[16 : 13];
  assign _zz_A_25 = ($signed(_zz__zz_A_25) + $signed(_zz__zz_A_25_1));
  assign _zz_A_26 = (_zz_when_LeakyRelu_l101_12 >>> 17);
  assign _zz_when_LeakyRelu_l101_12 = mul_6_P;
  assign when_LeakyRelu_l100_6 = _zz_when_LeakyRelu_l100_27[15];
  assign when_LeakyRelu_l101_6 = ($signed(_zz_when_LeakyRelu_l101_13) == $signed(_zz_when_LeakyRelu_l101_6_1));
  assign when_LeakyRelu_l104_6 = _zz_when_LeakyRelu_l101_12[16];
  assign when_LeakyRelu_l110_6 = (4'b1000 < _zz_when_LeakyRelu_l101_13);
  assign when_LeakyRelu_l103_6 = _zz_when_LeakyRelu_l101_12[17];
  assign when_LeakyRelu_l127_6 = _zz_when_LeakyRelu_l100_27_regNext[15];
  assign when_LeakyRelu_l131_96 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_96 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_97 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_97 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_98 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_98 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_99 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_99 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_100 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_100 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_101 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_101 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_102 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_102 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_103 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_103 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_104 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_104 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_105 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_105 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_106 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_106 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_107 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_107 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_108 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_108 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_109 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_109 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_110 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_110 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_111 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_111 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_6_1 = addSub_13_S;
  assign when_LeakyRelu_l155_6 = _zz_dataOut_6_1[15];
  assign when_LeakyRelu_l157_6 = ($signed(_zz_when_LeakyRelu_l157_6) < $signed(_zz_dataOut_6_1));
  assign dataOut_6 = _zz_dataOut_6;
  assign addSub_14_A = {8'h0,dataIn_7};
  assign _zz_when_LeakyRelu_l100_28 = addSub_14_S;
  assign _zz_when_LeakyRelu_l101_15 = _zz_when_LeakyRelu_l101_14[16 : 13];
  assign _zz_A_29 = ($signed(_zz__zz_A_29) + $signed(_zz__zz_A_29_1));
  assign _zz_A_30 = (_zz_when_LeakyRelu_l101_14 >>> 17);
  assign _zz_when_LeakyRelu_l101_14 = mul_7_P;
  assign when_LeakyRelu_l100_7 = _zz_when_LeakyRelu_l100_31[15];
  assign when_LeakyRelu_l101_7 = ($signed(_zz_when_LeakyRelu_l101_15) == $signed(_zz_when_LeakyRelu_l101_7_1));
  assign when_LeakyRelu_l104_7 = _zz_when_LeakyRelu_l101_14[16];
  assign when_LeakyRelu_l110_7 = (4'b1000 < _zz_when_LeakyRelu_l101_15);
  assign when_LeakyRelu_l103_7 = _zz_when_LeakyRelu_l101_14[17];
  assign when_LeakyRelu_l127_7 = _zz_when_LeakyRelu_l100_31_regNext[15];
  assign when_LeakyRelu_l131_112 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_112 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_113 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_113 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_114 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_114 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_115 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_115 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_116 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_116 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_117 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_117 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_118 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_118 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_119 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_119 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_120 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_120 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_121 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_121 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_122 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_122 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_123 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_123 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_124 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_124 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_125 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_125 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_126 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_126 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_127 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_127 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_7_1 = addSub_15_S;
  assign when_LeakyRelu_l155_7 = _zz_dataOut_7_1[15];
  assign when_LeakyRelu_l157_7 = ($signed(_zz_when_LeakyRelu_l157_7) < $signed(_zz_dataOut_7_1));
  assign dataOut_7 = _zz_dataOut_7;
  assign addSub_16_A = {8'h0,dataIn_8};
  assign _zz_when_LeakyRelu_l100_32 = addSub_16_S;
  assign _zz_when_LeakyRelu_l101_17 = _zz_when_LeakyRelu_l101_16[16 : 13];
  assign _zz_A_33 = ($signed(_zz__zz_A_33) + $signed(_zz__zz_A_33_1));
  assign _zz_A_34 = (_zz_when_LeakyRelu_l101_16 >>> 17);
  assign _zz_when_LeakyRelu_l101_16 = mul_8_P;
  assign when_LeakyRelu_l100_8 = _zz_when_LeakyRelu_l100_35[15];
  assign when_LeakyRelu_l101_8 = ($signed(_zz_when_LeakyRelu_l101_17) == $signed(_zz_when_LeakyRelu_l101_8_1));
  assign when_LeakyRelu_l104_8 = _zz_when_LeakyRelu_l101_16[16];
  assign when_LeakyRelu_l110_8 = (4'b1000 < _zz_when_LeakyRelu_l101_17);
  assign when_LeakyRelu_l103_8 = _zz_when_LeakyRelu_l101_16[17];
  assign when_LeakyRelu_l127_8 = _zz_when_LeakyRelu_l100_35_regNext[15];
  assign when_LeakyRelu_l131_128 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_128 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_129 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_129 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_130 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_130 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_131 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_131 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_132 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_132 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_133 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_133 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_134 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_134 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_135 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_135 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_136 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_136 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_137 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_137 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_138 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_138 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_139 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_139 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_140 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_140 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_141 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_141 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_142 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_142 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_143 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_143 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_8_1 = addSub_17_S;
  assign when_LeakyRelu_l155_8 = _zz_dataOut_8_1[15];
  assign when_LeakyRelu_l157_8 = ($signed(_zz_when_LeakyRelu_l157_8) < $signed(_zz_dataOut_8_1));
  assign dataOut_8 = _zz_dataOut_8;
  assign addSub_18_A = {8'h0,dataIn_9};
  assign _zz_when_LeakyRelu_l100_36 = addSub_18_S;
  assign _zz_when_LeakyRelu_l101_19 = _zz_when_LeakyRelu_l101_18[16 : 13];
  assign _zz_A_37 = ($signed(_zz__zz_A_37) + $signed(_zz__zz_A_37_1));
  assign _zz_A_38 = (_zz_when_LeakyRelu_l101_18 >>> 17);
  assign _zz_when_LeakyRelu_l101_18 = mul_9_P;
  assign when_LeakyRelu_l100_9 = _zz_when_LeakyRelu_l100_39[15];
  assign when_LeakyRelu_l101_9 = ($signed(_zz_when_LeakyRelu_l101_19) == $signed(_zz_when_LeakyRelu_l101_9_1));
  assign when_LeakyRelu_l104_9 = _zz_when_LeakyRelu_l101_18[16];
  assign when_LeakyRelu_l110_9 = (4'b1000 < _zz_when_LeakyRelu_l101_19);
  assign when_LeakyRelu_l103_9 = _zz_when_LeakyRelu_l101_18[17];
  assign when_LeakyRelu_l127_9 = _zz_when_LeakyRelu_l100_39_regNext[15];
  assign when_LeakyRelu_l131_144 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_144 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_145 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_145 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_146 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_146 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_147 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_147 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_148 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_148 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_149 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_149 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_150 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_150 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_151 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_151 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_152 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_152 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_153 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_153 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_154 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_154 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_155 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_155 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_156 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_156 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_157 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_157 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_158 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_158 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_159 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_159 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_9_1 = addSub_19_S;
  assign when_LeakyRelu_l155_9 = _zz_dataOut_9_1[15];
  assign when_LeakyRelu_l157_9 = ($signed(_zz_when_LeakyRelu_l157_9) < $signed(_zz_dataOut_9_1));
  assign dataOut_9 = _zz_dataOut_9;
  assign addSub_20_A = {8'h0,dataIn_10};
  assign _zz_when_LeakyRelu_l100_40 = addSub_20_S;
  assign _zz_when_LeakyRelu_l101_21 = _zz_when_LeakyRelu_l101_20[16 : 13];
  assign _zz_A_41 = ($signed(_zz__zz_A_41) + $signed(_zz__zz_A_41_1));
  assign _zz_A_42 = (_zz_when_LeakyRelu_l101_20 >>> 17);
  assign _zz_when_LeakyRelu_l101_20 = mul_10_P;
  assign when_LeakyRelu_l100_10 = _zz_when_LeakyRelu_l100_43[15];
  assign when_LeakyRelu_l101_10 = ($signed(_zz_when_LeakyRelu_l101_21) == $signed(_zz_when_LeakyRelu_l101_10_1));
  assign when_LeakyRelu_l104_10 = _zz_when_LeakyRelu_l101_20[16];
  assign when_LeakyRelu_l110_10 = (4'b1000 < _zz_when_LeakyRelu_l101_21);
  assign when_LeakyRelu_l103_10 = _zz_when_LeakyRelu_l101_20[17];
  assign when_LeakyRelu_l127_10 = _zz_when_LeakyRelu_l100_43_regNext[15];
  assign when_LeakyRelu_l131_160 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_160 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_161 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_161 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_162 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_162 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_163 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_163 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_164 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_164 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_165 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_165 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_166 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_166 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_167 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_167 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_168 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_168 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_169 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_169 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_170 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_170 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_171 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_171 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_172 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_172 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_173 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_173 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_174 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_174 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_175 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_175 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_10_1 = addSub_21_S;
  assign when_LeakyRelu_l155_10 = _zz_dataOut_10_1[15];
  assign when_LeakyRelu_l157_10 = ($signed(_zz_when_LeakyRelu_l157_10) < $signed(_zz_dataOut_10_1));
  assign dataOut_10 = _zz_dataOut_10;
  assign addSub_22_A = {8'h0,dataIn_11};
  assign _zz_when_LeakyRelu_l100_44 = addSub_22_S;
  assign _zz_when_LeakyRelu_l101_23 = _zz_when_LeakyRelu_l101_22[16 : 13];
  assign _zz_A_45 = ($signed(_zz__zz_A_45) + $signed(_zz__zz_A_45_1));
  assign _zz_A_46 = (_zz_when_LeakyRelu_l101_22 >>> 17);
  assign _zz_when_LeakyRelu_l101_22 = mul_11_P;
  assign when_LeakyRelu_l100_11 = _zz_when_LeakyRelu_l100_47[15];
  assign when_LeakyRelu_l101_11 = ($signed(_zz_when_LeakyRelu_l101_23) == $signed(_zz_when_LeakyRelu_l101_11_1));
  assign when_LeakyRelu_l104_11 = _zz_when_LeakyRelu_l101_22[16];
  assign when_LeakyRelu_l110_11 = (4'b1000 < _zz_when_LeakyRelu_l101_23);
  assign when_LeakyRelu_l103_11 = _zz_when_LeakyRelu_l101_22[17];
  assign when_LeakyRelu_l127_11 = _zz_when_LeakyRelu_l100_47_regNext[15];
  assign when_LeakyRelu_l131_176 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_176 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_177 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_177 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_178 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_178 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_179 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_179 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_180 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_180 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_181 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_181 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_182 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_182 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_183 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_183 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_184 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_184 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_185 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_185 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_186 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_186 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_187 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_187 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_188 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_188 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_189 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_189 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_190 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_190 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_191 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_191 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_11_1 = addSub_23_S;
  assign when_LeakyRelu_l155_11 = _zz_dataOut_11_1[15];
  assign when_LeakyRelu_l157_11 = ($signed(_zz_when_LeakyRelu_l157_11) < $signed(_zz_dataOut_11_1));
  assign dataOut_11 = _zz_dataOut_11;
  assign addSub_24_A = {8'h0,dataIn_12};
  assign _zz_when_LeakyRelu_l100_48 = addSub_24_S;
  assign _zz_when_LeakyRelu_l101_25 = _zz_when_LeakyRelu_l101_24[16 : 13];
  assign _zz_A_49 = ($signed(_zz__zz_A_49) + $signed(_zz__zz_A_49_1));
  assign _zz_A_50 = (_zz_when_LeakyRelu_l101_24 >>> 17);
  assign _zz_when_LeakyRelu_l101_24 = mul_12_P;
  assign when_LeakyRelu_l100_12 = _zz_when_LeakyRelu_l100_51[15];
  assign when_LeakyRelu_l101_12 = ($signed(_zz_when_LeakyRelu_l101_25) == $signed(_zz_when_LeakyRelu_l101_12_1));
  assign when_LeakyRelu_l104_12 = _zz_when_LeakyRelu_l101_24[16];
  assign when_LeakyRelu_l110_12 = (4'b1000 < _zz_when_LeakyRelu_l101_25);
  assign when_LeakyRelu_l103_12 = _zz_when_LeakyRelu_l101_24[17];
  assign when_LeakyRelu_l127_12 = _zz_when_LeakyRelu_l100_51_regNext[15];
  assign when_LeakyRelu_l131_192 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_192 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_193 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_193 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_194 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_194 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_195 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_195 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_196 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_196 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_197 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_197 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_198 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_198 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_199 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_199 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_200 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_200 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_201 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_201 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_202 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_202 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_203 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_203 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_204 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_204 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_205 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_205 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_206 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_206 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_207 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_207 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_12_1 = addSub_25_S;
  assign when_LeakyRelu_l155_12 = _zz_dataOut_12_1[15];
  assign when_LeakyRelu_l157_12 = ($signed(_zz_when_LeakyRelu_l157_12) < $signed(_zz_dataOut_12_1));
  assign dataOut_12 = _zz_dataOut_12;
  assign addSub_26_A = {8'h0,dataIn_13};
  assign _zz_when_LeakyRelu_l100_52 = addSub_26_S;
  assign _zz_when_LeakyRelu_l101_27 = _zz_when_LeakyRelu_l101_26[16 : 13];
  assign _zz_A_53 = ($signed(_zz__zz_A_53) + $signed(_zz__zz_A_53_1));
  assign _zz_A_54 = (_zz_when_LeakyRelu_l101_26 >>> 17);
  assign _zz_when_LeakyRelu_l101_26 = mul_13_P;
  assign when_LeakyRelu_l100_13 = _zz_when_LeakyRelu_l100_55[15];
  assign when_LeakyRelu_l101_13 = ($signed(_zz_when_LeakyRelu_l101_27) == $signed(_zz_when_LeakyRelu_l101_13_1));
  assign when_LeakyRelu_l104_13 = _zz_when_LeakyRelu_l101_26[16];
  assign when_LeakyRelu_l110_13 = (4'b1000 < _zz_when_LeakyRelu_l101_27);
  assign when_LeakyRelu_l103_13 = _zz_when_LeakyRelu_l101_26[17];
  assign when_LeakyRelu_l127_13 = _zz_when_LeakyRelu_l100_55_regNext[15];
  assign when_LeakyRelu_l131_208 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_208 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_209 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_209 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_210 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_210 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_211 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_211 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_212 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_212 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_213 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_213 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_214 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_214 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_215 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_215 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_216 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_216 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_217 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_217 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_218 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_218 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_219 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_219 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_220 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_220 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_221 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_221 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_222 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_222 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_223 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_223 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_13_1 = addSub_27_S;
  assign when_LeakyRelu_l155_13 = _zz_dataOut_13_1[15];
  assign when_LeakyRelu_l157_13 = ($signed(_zz_when_LeakyRelu_l157_13) < $signed(_zz_dataOut_13_1));
  assign dataOut_13 = _zz_dataOut_13;
  assign addSub_28_A = {8'h0,dataIn_14};
  assign _zz_when_LeakyRelu_l100_56 = addSub_28_S;
  assign _zz_when_LeakyRelu_l101_29 = _zz_when_LeakyRelu_l101_28[16 : 13];
  assign _zz_A_57 = ($signed(_zz__zz_A_57) + $signed(_zz__zz_A_57_1));
  assign _zz_A_58 = (_zz_when_LeakyRelu_l101_28 >>> 17);
  assign _zz_when_LeakyRelu_l101_28 = mul_14_P;
  assign when_LeakyRelu_l100_14 = _zz_when_LeakyRelu_l100_59[15];
  assign when_LeakyRelu_l101_14 = ($signed(_zz_when_LeakyRelu_l101_29) == $signed(_zz_when_LeakyRelu_l101_14_1));
  assign when_LeakyRelu_l104_14 = _zz_when_LeakyRelu_l101_28[16];
  assign when_LeakyRelu_l110_14 = (4'b1000 < _zz_when_LeakyRelu_l101_29);
  assign when_LeakyRelu_l103_14 = _zz_when_LeakyRelu_l101_28[17];
  assign when_LeakyRelu_l127_14 = _zz_when_LeakyRelu_l100_59_regNext[15];
  assign when_LeakyRelu_l131_224 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_224 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_225 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_225 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_226 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_226 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_227 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_227 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_228 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_228 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_229 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_229 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_230 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_230 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_231 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_231 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_232 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_232 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_233 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_233 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_234 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_234 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_235 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_235 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_236 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_236 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_237 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_237 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_238 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_238 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_239 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_239 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_14_1 = addSub_29_S;
  assign when_LeakyRelu_l155_14 = _zz_dataOut_14_1[15];
  assign when_LeakyRelu_l157_14 = ($signed(_zz_when_LeakyRelu_l157_14) < $signed(_zz_dataOut_14_1));
  assign dataOut_14 = _zz_dataOut_14;
  assign addSub_30_A = {8'h0,dataIn_15};
  assign _zz_when_LeakyRelu_l100_60 = addSub_30_S;
  assign _zz_when_LeakyRelu_l101_31 = _zz_when_LeakyRelu_l101_30[16 : 13];
  assign _zz_A_61 = ($signed(_zz__zz_A_61) + $signed(_zz__zz_A_61_1));
  assign _zz_A_62 = (_zz_when_LeakyRelu_l101_30 >>> 17);
  assign _zz_when_LeakyRelu_l101_30 = mul_15_P;
  assign when_LeakyRelu_l100_15 = _zz_when_LeakyRelu_l100_63[15];
  assign when_LeakyRelu_l101_15 = ($signed(_zz_when_LeakyRelu_l101_31) == $signed(_zz_when_LeakyRelu_l101_15_1));
  assign when_LeakyRelu_l104_15 = _zz_when_LeakyRelu_l101_30[16];
  assign when_LeakyRelu_l110_15 = (4'b1000 < _zz_when_LeakyRelu_l101_31);
  assign when_LeakyRelu_l103_15 = _zz_when_LeakyRelu_l101_30[17];
  assign when_LeakyRelu_l127_15 = _zz_when_LeakyRelu_l100_63_regNext[15];
  assign when_LeakyRelu_l131_240 = (amendReg[31 : 30] == 2'b01);
  assign when_LeakyRelu_l133_240 = (amendReg[31 : 30] == 2'b10);
  assign when_LeakyRelu_l131_241 = (amendReg[29 : 28] == 2'b01);
  assign when_LeakyRelu_l133_241 = (amendReg[29 : 28] == 2'b10);
  assign when_LeakyRelu_l131_242 = (amendReg[27 : 26] == 2'b01);
  assign when_LeakyRelu_l133_242 = (amendReg[27 : 26] == 2'b10);
  assign when_LeakyRelu_l131_243 = (amendReg[25 : 24] == 2'b01);
  assign when_LeakyRelu_l133_243 = (amendReg[25 : 24] == 2'b10);
  assign when_LeakyRelu_l131_244 = (amendReg[23 : 22] == 2'b01);
  assign when_LeakyRelu_l133_244 = (amendReg[23 : 22] == 2'b10);
  assign when_LeakyRelu_l131_245 = (amendReg[21 : 20] == 2'b01);
  assign when_LeakyRelu_l133_245 = (amendReg[21 : 20] == 2'b10);
  assign when_LeakyRelu_l131_246 = (amendReg[19 : 18] == 2'b01);
  assign when_LeakyRelu_l133_246 = (amendReg[19 : 18] == 2'b10);
  assign when_LeakyRelu_l131_247 = (amendReg[17 : 16] == 2'b01);
  assign when_LeakyRelu_l133_247 = (amendReg[17 : 16] == 2'b10);
  assign when_LeakyRelu_l131_248 = (amendReg[15 : 14] == 2'b01);
  assign when_LeakyRelu_l133_248 = (amendReg[15 : 14] == 2'b10);
  assign when_LeakyRelu_l131_249 = (amendReg[13 : 12] == 2'b01);
  assign when_LeakyRelu_l133_249 = (amendReg[13 : 12] == 2'b10);
  assign when_LeakyRelu_l131_250 = (amendReg[11 : 10] == 2'b01);
  assign when_LeakyRelu_l133_250 = (amendReg[11 : 10] == 2'b10);
  assign when_LeakyRelu_l131_251 = (amendReg[9 : 8] == 2'b01);
  assign when_LeakyRelu_l133_251 = (amendReg[9 : 8] == 2'b10);
  assign when_LeakyRelu_l131_252 = (amendReg[7 : 6] == 2'b01);
  assign when_LeakyRelu_l133_252 = (amendReg[7 : 6] == 2'b10);
  assign when_LeakyRelu_l131_253 = (amendReg[5 : 4] == 2'b01);
  assign when_LeakyRelu_l133_253 = (amendReg[5 : 4] == 2'b10);
  assign when_LeakyRelu_l131_254 = (amendReg[3 : 2] == 2'b01);
  assign when_LeakyRelu_l133_254 = (amendReg[3 : 2] == 2'b10);
  assign when_LeakyRelu_l131_255 = (amendReg[1 : 0] == 2'b01);
  assign when_LeakyRelu_l133_255 = (amendReg[1 : 0] == 2'b10);
  assign _zz_dataOut_15_1 = addSub_31_S;
  assign when_LeakyRelu_l155_15 = _zz_dataOut_15_1[15];
  assign when_LeakyRelu_l157_15 = ($signed(_zz_when_LeakyRelu_l157_15) < $signed(_zz_dataOut_15_1));
  assign dataOut_15 = _zz_dataOut_15;
  always @(posedge clk) begin
    _zz_when_LeakyRelu_l100_1 <= _zz_when_LeakyRelu_l100;
    _zz_when_LeakyRelu_l100_2 <= _zz_when_LeakyRelu_l100_1;
    _zz_when_LeakyRelu_l100_3 <= _zz_when_LeakyRelu_l100_2;
    if(when_LeakyRelu_l100) begin
      if(when_LeakyRelu_l101) begin
        _zz_A <= {{1{_zz_A_2[14]}}, _zz_A_2};
      end else begin
        if(when_LeakyRelu_l103) begin
          if(when_LeakyRelu_l104) begin
            _zz_A <= {{1{_zz_A_1[14]}}, _zz_A_1};
          end else begin
            _zz_A <= {{1{_zz_A_2[14]}}, _zz_A_2};
          end
        end else begin
          if(when_LeakyRelu_l110) begin
            _zz_A <= {{1{_zz_A_1[14]}}, _zz_A_1};
          end else begin
            _zz_A <= {{1{_zz_A_2[14]}}, _zz_A_2};
          end
        end
      end
    end else begin
      _zz_A <= _zz_when_LeakyRelu_l100_3;
    end
    _zz_when_LeakyRelu_l100_3_regNext <= _zz_when_LeakyRelu_l100_3;
    if(when_LeakyRelu_l127) begin
      case(_zz_when_LeakyRelu_l100_3_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3));
          end else begin
            if(when_LeakyRelu_l133) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_1));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_1) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_2));
          end else begin
            if(when_LeakyRelu_l133_1) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_3));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_2) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_4));
          end else begin
            if(when_LeakyRelu_l133_2) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_5));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_3) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_6));
          end else begin
            if(when_LeakyRelu_l133_3) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_7));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_4) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_8));
          end else begin
            if(when_LeakyRelu_l133_4) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_9));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_5) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_10));
          end else begin
            if(when_LeakyRelu_l133_5) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_11));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_6) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_12));
          end else begin
            if(when_LeakyRelu_l133_6) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_13));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_7) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_14));
          end else begin
            if(when_LeakyRelu_l133_7) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_15));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_8) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_16));
          end else begin
            if(when_LeakyRelu_l133_8) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_17));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_9) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_18));
          end else begin
            if(when_LeakyRelu_l133_9) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_19));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_10) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_20));
          end else begin
            if(when_LeakyRelu_l133_10) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_21));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_11) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_22));
          end else begin
            if(when_LeakyRelu_l133_11) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_23));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_12) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_24));
          end else begin
            if(when_LeakyRelu_l133_12) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_25));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_13) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_26));
          end else begin
            if(when_LeakyRelu_l133_13) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_27));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_14) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_28));
          end else begin
            if(when_LeakyRelu_l133_14) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_29));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_15) begin
            _zz_A_3 <= ($signed(_zz_A) + $signed(_zz__zz_A_3_30));
          end else begin
            if(when_LeakyRelu_l133_15) begin
              _zz_A_3 <= ($signed(_zz_A) - $signed(_zz__zz_A_3_31));
            end else begin
              _zz_A_3 <= _zz_A;
            end
          end
        end
        default : begin
          _zz_A_3 <= _zz_A;
        end
      endcase
    end else begin
      _zz_A_3 <= _zz_A;
    end
    if(when_LeakyRelu_l155) begin
      _zz_dataOut_0 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157) begin
        _zz_dataOut_0 <= 8'hff;
      end else begin
        _zz_dataOut_0 <= _zz__zz_dataOut_0[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_5 <= _zz_when_LeakyRelu_l100_4;
    _zz_when_LeakyRelu_l100_6 <= _zz_when_LeakyRelu_l100_5;
    _zz_when_LeakyRelu_l100_7 <= _zz_when_LeakyRelu_l100_6;
    if(when_LeakyRelu_l100_1) begin
      if(when_LeakyRelu_l101_1) begin
        _zz_A_4 <= {{1{_zz_A_6[14]}}, _zz_A_6};
      end else begin
        if(when_LeakyRelu_l103_1) begin
          if(when_LeakyRelu_l104_1) begin
            _zz_A_4 <= {{1{_zz_A_5[14]}}, _zz_A_5};
          end else begin
            _zz_A_4 <= {{1{_zz_A_6[14]}}, _zz_A_6};
          end
        end else begin
          if(when_LeakyRelu_l110_1) begin
            _zz_A_4 <= {{1{_zz_A_5[14]}}, _zz_A_5};
          end else begin
            _zz_A_4 <= {{1{_zz_A_6[14]}}, _zz_A_6};
          end
        end
      end
    end else begin
      _zz_A_4 <= _zz_when_LeakyRelu_l100_7;
    end
    _zz_when_LeakyRelu_l100_7_regNext <= _zz_when_LeakyRelu_l100_7;
    if(when_LeakyRelu_l127_1) begin
      case(_zz_when_LeakyRelu_l100_7_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_16) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7));
          end else begin
            if(when_LeakyRelu_l133_16) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_1));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_17) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_2));
          end else begin
            if(when_LeakyRelu_l133_17) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_3));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_18) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_4));
          end else begin
            if(when_LeakyRelu_l133_18) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_5));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_19) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_6));
          end else begin
            if(when_LeakyRelu_l133_19) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_7));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_20) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_8));
          end else begin
            if(when_LeakyRelu_l133_20) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_9));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_21) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_10));
          end else begin
            if(when_LeakyRelu_l133_21) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_11));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_22) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_12));
          end else begin
            if(when_LeakyRelu_l133_22) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_13));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_23) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_14));
          end else begin
            if(when_LeakyRelu_l133_23) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_15));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_24) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_16));
          end else begin
            if(when_LeakyRelu_l133_24) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_17));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_25) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_18));
          end else begin
            if(when_LeakyRelu_l133_25) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_19));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_26) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_20));
          end else begin
            if(when_LeakyRelu_l133_26) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_21));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_27) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_22));
          end else begin
            if(when_LeakyRelu_l133_27) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_23));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_28) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_24));
          end else begin
            if(when_LeakyRelu_l133_28) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_25));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_29) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_26));
          end else begin
            if(when_LeakyRelu_l133_29) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_27));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_30) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_28));
          end else begin
            if(when_LeakyRelu_l133_30) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_29));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_31) begin
            _zz_A_7 <= ($signed(_zz_A_4) + $signed(_zz__zz_A_7_30));
          end else begin
            if(when_LeakyRelu_l133_31) begin
              _zz_A_7 <= ($signed(_zz_A_4) - $signed(_zz__zz_A_7_31));
            end else begin
              _zz_A_7 <= _zz_A_4;
            end
          end
        end
        default : begin
          _zz_A_7 <= _zz_A_4;
        end
      endcase
    end else begin
      _zz_A_7 <= _zz_A_4;
    end
    if(when_LeakyRelu_l155_1) begin
      _zz_dataOut_1 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_1) begin
        _zz_dataOut_1 <= 8'hff;
      end else begin
        _zz_dataOut_1 <= _zz__zz_dataOut_1[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_9 <= _zz_when_LeakyRelu_l100_8;
    _zz_when_LeakyRelu_l100_10 <= _zz_when_LeakyRelu_l100_9;
    _zz_when_LeakyRelu_l100_11 <= _zz_when_LeakyRelu_l100_10;
    if(when_LeakyRelu_l100_2) begin
      if(when_LeakyRelu_l101_2) begin
        _zz_A_8 <= {{1{_zz_A_10[14]}}, _zz_A_10};
      end else begin
        if(when_LeakyRelu_l103_2) begin
          if(when_LeakyRelu_l104_2) begin
            _zz_A_8 <= {{1{_zz_A_9[14]}}, _zz_A_9};
          end else begin
            _zz_A_8 <= {{1{_zz_A_10[14]}}, _zz_A_10};
          end
        end else begin
          if(when_LeakyRelu_l110_2) begin
            _zz_A_8 <= {{1{_zz_A_9[14]}}, _zz_A_9};
          end else begin
            _zz_A_8 <= {{1{_zz_A_10[14]}}, _zz_A_10};
          end
        end
      end
    end else begin
      _zz_A_8 <= _zz_when_LeakyRelu_l100_11;
    end
    _zz_when_LeakyRelu_l100_11_regNext <= _zz_when_LeakyRelu_l100_11;
    if(when_LeakyRelu_l127_2) begin
      case(_zz_when_LeakyRelu_l100_11_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_32) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11));
          end else begin
            if(when_LeakyRelu_l133_32) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_1));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_33) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_2));
          end else begin
            if(when_LeakyRelu_l133_33) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_3));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_34) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_4));
          end else begin
            if(when_LeakyRelu_l133_34) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_5));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_35) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_6));
          end else begin
            if(when_LeakyRelu_l133_35) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_7));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_36) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_8));
          end else begin
            if(when_LeakyRelu_l133_36) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_9));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_37) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_10));
          end else begin
            if(when_LeakyRelu_l133_37) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_11));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_38) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_12));
          end else begin
            if(when_LeakyRelu_l133_38) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_13));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_39) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_14));
          end else begin
            if(when_LeakyRelu_l133_39) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_15));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_40) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_16));
          end else begin
            if(when_LeakyRelu_l133_40) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_17));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_41) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_18));
          end else begin
            if(when_LeakyRelu_l133_41) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_19));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_42) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_20));
          end else begin
            if(when_LeakyRelu_l133_42) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_21));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_43) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_22));
          end else begin
            if(when_LeakyRelu_l133_43) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_23));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_44) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_24));
          end else begin
            if(when_LeakyRelu_l133_44) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_25));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_45) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_26));
          end else begin
            if(when_LeakyRelu_l133_45) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_27));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_46) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_28));
          end else begin
            if(when_LeakyRelu_l133_46) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_29));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_47) begin
            _zz_A_11 <= ($signed(_zz_A_8) + $signed(_zz__zz_A_11_30));
          end else begin
            if(when_LeakyRelu_l133_47) begin
              _zz_A_11 <= ($signed(_zz_A_8) - $signed(_zz__zz_A_11_31));
            end else begin
              _zz_A_11 <= _zz_A_8;
            end
          end
        end
        default : begin
          _zz_A_11 <= _zz_A_8;
        end
      endcase
    end else begin
      _zz_A_11 <= _zz_A_8;
    end
    if(when_LeakyRelu_l155_2) begin
      _zz_dataOut_2 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_2) begin
        _zz_dataOut_2 <= 8'hff;
      end else begin
        _zz_dataOut_2 <= _zz__zz_dataOut_2[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_13 <= _zz_when_LeakyRelu_l100_12;
    _zz_when_LeakyRelu_l100_14 <= _zz_when_LeakyRelu_l100_13;
    _zz_when_LeakyRelu_l100_15 <= _zz_when_LeakyRelu_l100_14;
    if(when_LeakyRelu_l100_3) begin
      if(when_LeakyRelu_l101_3) begin
        _zz_A_12 <= {{1{_zz_A_14[14]}}, _zz_A_14};
      end else begin
        if(when_LeakyRelu_l103_3) begin
          if(when_LeakyRelu_l104_3) begin
            _zz_A_12 <= {{1{_zz_A_13[14]}}, _zz_A_13};
          end else begin
            _zz_A_12 <= {{1{_zz_A_14[14]}}, _zz_A_14};
          end
        end else begin
          if(when_LeakyRelu_l110_3) begin
            _zz_A_12 <= {{1{_zz_A_13[14]}}, _zz_A_13};
          end else begin
            _zz_A_12 <= {{1{_zz_A_14[14]}}, _zz_A_14};
          end
        end
      end
    end else begin
      _zz_A_12 <= _zz_when_LeakyRelu_l100_15;
    end
    _zz_when_LeakyRelu_l100_15_regNext <= _zz_when_LeakyRelu_l100_15;
    if(when_LeakyRelu_l127_3) begin
      case(_zz_when_LeakyRelu_l100_15_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_48) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15));
          end else begin
            if(when_LeakyRelu_l133_48) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_1));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_49) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_2));
          end else begin
            if(when_LeakyRelu_l133_49) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_3));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_50) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_4));
          end else begin
            if(when_LeakyRelu_l133_50) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_5));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_51) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_6));
          end else begin
            if(when_LeakyRelu_l133_51) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_7));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_52) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_8));
          end else begin
            if(when_LeakyRelu_l133_52) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_9));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_53) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_10));
          end else begin
            if(when_LeakyRelu_l133_53) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_11));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_54) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_12));
          end else begin
            if(when_LeakyRelu_l133_54) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_13));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_55) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_14));
          end else begin
            if(when_LeakyRelu_l133_55) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_15));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_56) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_16));
          end else begin
            if(when_LeakyRelu_l133_56) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_17));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_57) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_18));
          end else begin
            if(when_LeakyRelu_l133_57) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_19));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_58) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_20));
          end else begin
            if(when_LeakyRelu_l133_58) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_21));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_59) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_22));
          end else begin
            if(when_LeakyRelu_l133_59) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_23));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_60) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_24));
          end else begin
            if(when_LeakyRelu_l133_60) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_25));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_61) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_26));
          end else begin
            if(when_LeakyRelu_l133_61) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_27));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_62) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_28));
          end else begin
            if(when_LeakyRelu_l133_62) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_29));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_63) begin
            _zz_A_15 <= ($signed(_zz_A_12) + $signed(_zz__zz_A_15_30));
          end else begin
            if(when_LeakyRelu_l133_63) begin
              _zz_A_15 <= ($signed(_zz_A_12) - $signed(_zz__zz_A_15_31));
            end else begin
              _zz_A_15 <= _zz_A_12;
            end
          end
        end
        default : begin
          _zz_A_15 <= _zz_A_12;
        end
      endcase
    end else begin
      _zz_A_15 <= _zz_A_12;
    end
    if(when_LeakyRelu_l155_3) begin
      _zz_dataOut_3 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_3) begin
        _zz_dataOut_3 <= 8'hff;
      end else begin
        _zz_dataOut_3 <= _zz__zz_dataOut_3[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_17 <= _zz_when_LeakyRelu_l100_16;
    _zz_when_LeakyRelu_l100_18 <= _zz_when_LeakyRelu_l100_17;
    _zz_when_LeakyRelu_l100_19 <= _zz_when_LeakyRelu_l100_18;
    if(when_LeakyRelu_l100_4) begin
      if(when_LeakyRelu_l101_4) begin
        _zz_A_16 <= {{1{_zz_A_18[14]}}, _zz_A_18};
      end else begin
        if(when_LeakyRelu_l103_4) begin
          if(when_LeakyRelu_l104_4) begin
            _zz_A_16 <= {{1{_zz_A_17[14]}}, _zz_A_17};
          end else begin
            _zz_A_16 <= {{1{_zz_A_18[14]}}, _zz_A_18};
          end
        end else begin
          if(when_LeakyRelu_l110_4) begin
            _zz_A_16 <= {{1{_zz_A_17[14]}}, _zz_A_17};
          end else begin
            _zz_A_16 <= {{1{_zz_A_18[14]}}, _zz_A_18};
          end
        end
      end
    end else begin
      _zz_A_16 <= _zz_when_LeakyRelu_l100_19;
    end
    _zz_when_LeakyRelu_l100_19_regNext <= _zz_when_LeakyRelu_l100_19;
    if(when_LeakyRelu_l127_4) begin
      case(_zz_when_LeakyRelu_l100_19_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_64) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19));
          end else begin
            if(when_LeakyRelu_l133_64) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_1));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_65) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_2));
          end else begin
            if(when_LeakyRelu_l133_65) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_3));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_66) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_4));
          end else begin
            if(when_LeakyRelu_l133_66) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_5));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_67) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_6));
          end else begin
            if(when_LeakyRelu_l133_67) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_7));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_68) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_8));
          end else begin
            if(when_LeakyRelu_l133_68) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_9));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_69) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_10));
          end else begin
            if(when_LeakyRelu_l133_69) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_11));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_70) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_12));
          end else begin
            if(when_LeakyRelu_l133_70) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_13));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_71) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_14));
          end else begin
            if(when_LeakyRelu_l133_71) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_15));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_72) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_16));
          end else begin
            if(when_LeakyRelu_l133_72) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_17));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_73) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_18));
          end else begin
            if(when_LeakyRelu_l133_73) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_19));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_74) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_20));
          end else begin
            if(when_LeakyRelu_l133_74) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_21));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_75) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_22));
          end else begin
            if(when_LeakyRelu_l133_75) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_23));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_76) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_24));
          end else begin
            if(when_LeakyRelu_l133_76) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_25));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_77) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_26));
          end else begin
            if(when_LeakyRelu_l133_77) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_27));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_78) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_28));
          end else begin
            if(when_LeakyRelu_l133_78) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_29));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_79) begin
            _zz_A_19 <= ($signed(_zz_A_16) + $signed(_zz__zz_A_19_30));
          end else begin
            if(when_LeakyRelu_l133_79) begin
              _zz_A_19 <= ($signed(_zz_A_16) - $signed(_zz__zz_A_19_31));
            end else begin
              _zz_A_19 <= _zz_A_16;
            end
          end
        end
        default : begin
          _zz_A_19 <= _zz_A_16;
        end
      endcase
    end else begin
      _zz_A_19 <= _zz_A_16;
    end
    if(when_LeakyRelu_l155_4) begin
      _zz_dataOut_4 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_4) begin
        _zz_dataOut_4 <= 8'hff;
      end else begin
        _zz_dataOut_4 <= _zz__zz_dataOut_4[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_21 <= _zz_when_LeakyRelu_l100_20;
    _zz_when_LeakyRelu_l100_22 <= _zz_when_LeakyRelu_l100_21;
    _zz_when_LeakyRelu_l100_23 <= _zz_when_LeakyRelu_l100_22;
    if(when_LeakyRelu_l100_5) begin
      if(when_LeakyRelu_l101_5) begin
        _zz_A_20 <= {{1{_zz_A_22[14]}}, _zz_A_22};
      end else begin
        if(when_LeakyRelu_l103_5) begin
          if(when_LeakyRelu_l104_5) begin
            _zz_A_20 <= {{1{_zz_A_21[14]}}, _zz_A_21};
          end else begin
            _zz_A_20 <= {{1{_zz_A_22[14]}}, _zz_A_22};
          end
        end else begin
          if(when_LeakyRelu_l110_5) begin
            _zz_A_20 <= {{1{_zz_A_21[14]}}, _zz_A_21};
          end else begin
            _zz_A_20 <= {{1{_zz_A_22[14]}}, _zz_A_22};
          end
        end
      end
    end else begin
      _zz_A_20 <= _zz_when_LeakyRelu_l100_23;
    end
    _zz_when_LeakyRelu_l100_23_regNext <= _zz_when_LeakyRelu_l100_23;
    if(when_LeakyRelu_l127_5) begin
      case(_zz_when_LeakyRelu_l100_23_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_80) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23));
          end else begin
            if(when_LeakyRelu_l133_80) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_1));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_81) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_2));
          end else begin
            if(when_LeakyRelu_l133_81) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_3));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_82) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_4));
          end else begin
            if(when_LeakyRelu_l133_82) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_5));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_83) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_6));
          end else begin
            if(when_LeakyRelu_l133_83) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_7));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_84) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_8));
          end else begin
            if(when_LeakyRelu_l133_84) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_9));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_85) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_10));
          end else begin
            if(when_LeakyRelu_l133_85) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_11));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_86) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_12));
          end else begin
            if(when_LeakyRelu_l133_86) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_13));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_87) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_14));
          end else begin
            if(when_LeakyRelu_l133_87) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_15));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_88) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_16));
          end else begin
            if(when_LeakyRelu_l133_88) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_17));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_89) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_18));
          end else begin
            if(when_LeakyRelu_l133_89) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_19));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_90) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_20));
          end else begin
            if(when_LeakyRelu_l133_90) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_21));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_91) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_22));
          end else begin
            if(when_LeakyRelu_l133_91) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_23));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_92) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_24));
          end else begin
            if(when_LeakyRelu_l133_92) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_25));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_93) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_26));
          end else begin
            if(when_LeakyRelu_l133_93) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_27));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_94) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_28));
          end else begin
            if(when_LeakyRelu_l133_94) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_29));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_95) begin
            _zz_A_23 <= ($signed(_zz_A_20) + $signed(_zz__zz_A_23_30));
          end else begin
            if(when_LeakyRelu_l133_95) begin
              _zz_A_23 <= ($signed(_zz_A_20) - $signed(_zz__zz_A_23_31));
            end else begin
              _zz_A_23 <= _zz_A_20;
            end
          end
        end
        default : begin
          _zz_A_23 <= _zz_A_20;
        end
      endcase
    end else begin
      _zz_A_23 <= _zz_A_20;
    end
    if(when_LeakyRelu_l155_5) begin
      _zz_dataOut_5 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_5) begin
        _zz_dataOut_5 <= 8'hff;
      end else begin
        _zz_dataOut_5 <= _zz__zz_dataOut_5[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_25 <= _zz_when_LeakyRelu_l100_24;
    _zz_when_LeakyRelu_l100_26 <= _zz_when_LeakyRelu_l100_25;
    _zz_when_LeakyRelu_l100_27 <= _zz_when_LeakyRelu_l100_26;
    if(when_LeakyRelu_l100_6) begin
      if(when_LeakyRelu_l101_6) begin
        _zz_A_24 <= {{1{_zz_A_26[14]}}, _zz_A_26};
      end else begin
        if(when_LeakyRelu_l103_6) begin
          if(when_LeakyRelu_l104_6) begin
            _zz_A_24 <= {{1{_zz_A_25[14]}}, _zz_A_25};
          end else begin
            _zz_A_24 <= {{1{_zz_A_26[14]}}, _zz_A_26};
          end
        end else begin
          if(when_LeakyRelu_l110_6) begin
            _zz_A_24 <= {{1{_zz_A_25[14]}}, _zz_A_25};
          end else begin
            _zz_A_24 <= {{1{_zz_A_26[14]}}, _zz_A_26};
          end
        end
      end
    end else begin
      _zz_A_24 <= _zz_when_LeakyRelu_l100_27;
    end
    _zz_when_LeakyRelu_l100_27_regNext <= _zz_when_LeakyRelu_l100_27;
    if(when_LeakyRelu_l127_6) begin
      case(_zz_when_LeakyRelu_l100_27_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_96) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27));
          end else begin
            if(when_LeakyRelu_l133_96) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_1));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_97) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_2));
          end else begin
            if(when_LeakyRelu_l133_97) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_3));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_98) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_4));
          end else begin
            if(when_LeakyRelu_l133_98) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_5));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_99) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_6));
          end else begin
            if(when_LeakyRelu_l133_99) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_7));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_100) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_8));
          end else begin
            if(when_LeakyRelu_l133_100) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_9));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_101) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_10));
          end else begin
            if(when_LeakyRelu_l133_101) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_11));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_102) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_12));
          end else begin
            if(when_LeakyRelu_l133_102) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_13));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_103) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_14));
          end else begin
            if(when_LeakyRelu_l133_103) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_15));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_104) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_16));
          end else begin
            if(when_LeakyRelu_l133_104) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_17));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_105) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_18));
          end else begin
            if(when_LeakyRelu_l133_105) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_19));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_106) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_20));
          end else begin
            if(when_LeakyRelu_l133_106) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_21));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_107) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_22));
          end else begin
            if(when_LeakyRelu_l133_107) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_23));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_108) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_24));
          end else begin
            if(when_LeakyRelu_l133_108) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_25));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_109) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_26));
          end else begin
            if(when_LeakyRelu_l133_109) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_27));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_110) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_28));
          end else begin
            if(when_LeakyRelu_l133_110) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_29));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_111) begin
            _zz_A_27 <= ($signed(_zz_A_24) + $signed(_zz__zz_A_27_30));
          end else begin
            if(when_LeakyRelu_l133_111) begin
              _zz_A_27 <= ($signed(_zz_A_24) - $signed(_zz__zz_A_27_31));
            end else begin
              _zz_A_27 <= _zz_A_24;
            end
          end
        end
        default : begin
          _zz_A_27 <= _zz_A_24;
        end
      endcase
    end else begin
      _zz_A_27 <= _zz_A_24;
    end
    if(when_LeakyRelu_l155_6) begin
      _zz_dataOut_6 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_6) begin
        _zz_dataOut_6 <= 8'hff;
      end else begin
        _zz_dataOut_6 <= _zz__zz_dataOut_6[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_29 <= _zz_when_LeakyRelu_l100_28;
    _zz_when_LeakyRelu_l100_30 <= _zz_when_LeakyRelu_l100_29;
    _zz_when_LeakyRelu_l100_31 <= _zz_when_LeakyRelu_l100_30;
    if(when_LeakyRelu_l100_7) begin
      if(when_LeakyRelu_l101_7) begin
        _zz_A_28 <= {{1{_zz_A_30[14]}}, _zz_A_30};
      end else begin
        if(when_LeakyRelu_l103_7) begin
          if(when_LeakyRelu_l104_7) begin
            _zz_A_28 <= {{1{_zz_A_29[14]}}, _zz_A_29};
          end else begin
            _zz_A_28 <= {{1{_zz_A_30[14]}}, _zz_A_30};
          end
        end else begin
          if(when_LeakyRelu_l110_7) begin
            _zz_A_28 <= {{1{_zz_A_29[14]}}, _zz_A_29};
          end else begin
            _zz_A_28 <= {{1{_zz_A_30[14]}}, _zz_A_30};
          end
        end
      end
    end else begin
      _zz_A_28 <= _zz_when_LeakyRelu_l100_31;
    end
    _zz_when_LeakyRelu_l100_31_regNext <= _zz_when_LeakyRelu_l100_31;
    if(when_LeakyRelu_l127_7) begin
      case(_zz_when_LeakyRelu_l100_31_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_112) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31));
          end else begin
            if(when_LeakyRelu_l133_112) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_1));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_113) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_2));
          end else begin
            if(when_LeakyRelu_l133_113) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_3));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_114) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_4));
          end else begin
            if(when_LeakyRelu_l133_114) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_5));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_115) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_6));
          end else begin
            if(when_LeakyRelu_l133_115) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_7));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_116) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_8));
          end else begin
            if(when_LeakyRelu_l133_116) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_9));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_117) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_10));
          end else begin
            if(when_LeakyRelu_l133_117) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_11));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_118) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_12));
          end else begin
            if(when_LeakyRelu_l133_118) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_13));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_119) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_14));
          end else begin
            if(when_LeakyRelu_l133_119) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_15));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_120) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_16));
          end else begin
            if(when_LeakyRelu_l133_120) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_17));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_121) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_18));
          end else begin
            if(when_LeakyRelu_l133_121) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_19));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_122) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_20));
          end else begin
            if(when_LeakyRelu_l133_122) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_21));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_123) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_22));
          end else begin
            if(when_LeakyRelu_l133_123) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_23));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_124) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_24));
          end else begin
            if(when_LeakyRelu_l133_124) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_25));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_125) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_26));
          end else begin
            if(when_LeakyRelu_l133_125) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_27));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_126) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_28));
          end else begin
            if(when_LeakyRelu_l133_126) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_29));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_127) begin
            _zz_A_31 <= ($signed(_zz_A_28) + $signed(_zz__zz_A_31_30));
          end else begin
            if(when_LeakyRelu_l133_127) begin
              _zz_A_31 <= ($signed(_zz_A_28) - $signed(_zz__zz_A_31_31));
            end else begin
              _zz_A_31 <= _zz_A_28;
            end
          end
        end
        default : begin
          _zz_A_31 <= _zz_A_28;
        end
      endcase
    end else begin
      _zz_A_31 <= _zz_A_28;
    end
    if(when_LeakyRelu_l155_7) begin
      _zz_dataOut_7 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_7) begin
        _zz_dataOut_7 <= 8'hff;
      end else begin
        _zz_dataOut_7 <= _zz__zz_dataOut_7[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_33 <= _zz_when_LeakyRelu_l100_32;
    _zz_when_LeakyRelu_l100_34 <= _zz_when_LeakyRelu_l100_33;
    _zz_when_LeakyRelu_l100_35 <= _zz_when_LeakyRelu_l100_34;
    if(when_LeakyRelu_l100_8) begin
      if(when_LeakyRelu_l101_8) begin
        _zz_A_32 <= {{1{_zz_A_34[14]}}, _zz_A_34};
      end else begin
        if(when_LeakyRelu_l103_8) begin
          if(when_LeakyRelu_l104_8) begin
            _zz_A_32 <= {{1{_zz_A_33[14]}}, _zz_A_33};
          end else begin
            _zz_A_32 <= {{1{_zz_A_34[14]}}, _zz_A_34};
          end
        end else begin
          if(when_LeakyRelu_l110_8) begin
            _zz_A_32 <= {{1{_zz_A_33[14]}}, _zz_A_33};
          end else begin
            _zz_A_32 <= {{1{_zz_A_34[14]}}, _zz_A_34};
          end
        end
      end
    end else begin
      _zz_A_32 <= _zz_when_LeakyRelu_l100_35;
    end
    _zz_when_LeakyRelu_l100_35_regNext <= _zz_when_LeakyRelu_l100_35;
    if(when_LeakyRelu_l127_8) begin
      case(_zz_when_LeakyRelu_l100_35_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_128) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35));
          end else begin
            if(when_LeakyRelu_l133_128) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_1));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_129) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_2));
          end else begin
            if(when_LeakyRelu_l133_129) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_3));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_130) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_4));
          end else begin
            if(when_LeakyRelu_l133_130) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_5));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_131) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_6));
          end else begin
            if(when_LeakyRelu_l133_131) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_7));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_132) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_8));
          end else begin
            if(when_LeakyRelu_l133_132) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_9));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_133) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_10));
          end else begin
            if(when_LeakyRelu_l133_133) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_11));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_134) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_12));
          end else begin
            if(when_LeakyRelu_l133_134) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_13));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_135) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_14));
          end else begin
            if(when_LeakyRelu_l133_135) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_15));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_136) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_16));
          end else begin
            if(when_LeakyRelu_l133_136) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_17));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_137) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_18));
          end else begin
            if(when_LeakyRelu_l133_137) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_19));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_138) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_20));
          end else begin
            if(when_LeakyRelu_l133_138) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_21));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_139) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_22));
          end else begin
            if(when_LeakyRelu_l133_139) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_23));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_140) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_24));
          end else begin
            if(when_LeakyRelu_l133_140) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_25));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_141) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_26));
          end else begin
            if(when_LeakyRelu_l133_141) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_27));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_142) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_28));
          end else begin
            if(when_LeakyRelu_l133_142) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_29));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_143) begin
            _zz_A_35 <= ($signed(_zz_A_32) + $signed(_zz__zz_A_35_30));
          end else begin
            if(when_LeakyRelu_l133_143) begin
              _zz_A_35 <= ($signed(_zz_A_32) - $signed(_zz__zz_A_35_31));
            end else begin
              _zz_A_35 <= _zz_A_32;
            end
          end
        end
        default : begin
          _zz_A_35 <= _zz_A_32;
        end
      endcase
    end else begin
      _zz_A_35 <= _zz_A_32;
    end
    if(when_LeakyRelu_l155_8) begin
      _zz_dataOut_8 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_8) begin
        _zz_dataOut_8 <= 8'hff;
      end else begin
        _zz_dataOut_8 <= _zz__zz_dataOut_8[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_37 <= _zz_when_LeakyRelu_l100_36;
    _zz_when_LeakyRelu_l100_38 <= _zz_when_LeakyRelu_l100_37;
    _zz_when_LeakyRelu_l100_39 <= _zz_when_LeakyRelu_l100_38;
    if(when_LeakyRelu_l100_9) begin
      if(when_LeakyRelu_l101_9) begin
        _zz_A_36 <= {{1{_zz_A_38[14]}}, _zz_A_38};
      end else begin
        if(when_LeakyRelu_l103_9) begin
          if(when_LeakyRelu_l104_9) begin
            _zz_A_36 <= {{1{_zz_A_37[14]}}, _zz_A_37};
          end else begin
            _zz_A_36 <= {{1{_zz_A_38[14]}}, _zz_A_38};
          end
        end else begin
          if(when_LeakyRelu_l110_9) begin
            _zz_A_36 <= {{1{_zz_A_37[14]}}, _zz_A_37};
          end else begin
            _zz_A_36 <= {{1{_zz_A_38[14]}}, _zz_A_38};
          end
        end
      end
    end else begin
      _zz_A_36 <= _zz_when_LeakyRelu_l100_39;
    end
    _zz_when_LeakyRelu_l100_39_regNext <= _zz_when_LeakyRelu_l100_39;
    if(when_LeakyRelu_l127_9) begin
      case(_zz_when_LeakyRelu_l100_39_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_144) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39));
          end else begin
            if(when_LeakyRelu_l133_144) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_1));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_145) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_2));
          end else begin
            if(when_LeakyRelu_l133_145) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_3));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_146) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_4));
          end else begin
            if(when_LeakyRelu_l133_146) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_5));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_147) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_6));
          end else begin
            if(when_LeakyRelu_l133_147) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_7));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_148) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_8));
          end else begin
            if(when_LeakyRelu_l133_148) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_9));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_149) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_10));
          end else begin
            if(when_LeakyRelu_l133_149) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_11));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_150) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_12));
          end else begin
            if(when_LeakyRelu_l133_150) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_13));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_151) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_14));
          end else begin
            if(when_LeakyRelu_l133_151) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_15));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_152) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_16));
          end else begin
            if(when_LeakyRelu_l133_152) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_17));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_153) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_18));
          end else begin
            if(when_LeakyRelu_l133_153) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_19));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_154) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_20));
          end else begin
            if(when_LeakyRelu_l133_154) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_21));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_155) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_22));
          end else begin
            if(when_LeakyRelu_l133_155) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_23));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_156) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_24));
          end else begin
            if(when_LeakyRelu_l133_156) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_25));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_157) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_26));
          end else begin
            if(when_LeakyRelu_l133_157) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_27));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_158) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_28));
          end else begin
            if(when_LeakyRelu_l133_158) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_29));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_159) begin
            _zz_A_39 <= ($signed(_zz_A_36) + $signed(_zz__zz_A_39_30));
          end else begin
            if(when_LeakyRelu_l133_159) begin
              _zz_A_39 <= ($signed(_zz_A_36) - $signed(_zz__zz_A_39_31));
            end else begin
              _zz_A_39 <= _zz_A_36;
            end
          end
        end
        default : begin
          _zz_A_39 <= _zz_A_36;
        end
      endcase
    end else begin
      _zz_A_39 <= _zz_A_36;
    end
    if(when_LeakyRelu_l155_9) begin
      _zz_dataOut_9 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_9) begin
        _zz_dataOut_9 <= 8'hff;
      end else begin
        _zz_dataOut_9 <= _zz__zz_dataOut_9[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_41 <= _zz_when_LeakyRelu_l100_40;
    _zz_when_LeakyRelu_l100_42 <= _zz_when_LeakyRelu_l100_41;
    _zz_when_LeakyRelu_l100_43 <= _zz_when_LeakyRelu_l100_42;
    if(when_LeakyRelu_l100_10) begin
      if(when_LeakyRelu_l101_10) begin
        _zz_A_40 <= {{1{_zz_A_42[14]}}, _zz_A_42};
      end else begin
        if(when_LeakyRelu_l103_10) begin
          if(when_LeakyRelu_l104_10) begin
            _zz_A_40 <= {{1{_zz_A_41[14]}}, _zz_A_41};
          end else begin
            _zz_A_40 <= {{1{_zz_A_42[14]}}, _zz_A_42};
          end
        end else begin
          if(when_LeakyRelu_l110_10) begin
            _zz_A_40 <= {{1{_zz_A_41[14]}}, _zz_A_41};
          end else begin
            _zz_A_40 <= {{1{_zz_A_42[14]}}, _zz_A_42};
          end
        end
      end
    end else begin
      _zz_A_40 <= _zz_when_LeakyRelu_l100_43;
    end
    _zz_when_LeakyRelu_l100_43_regNext <= _zz_when_LeakyRelu_l100_43;
    if(when_LeakyRelu_l127_10) begin
      case(_zz_when_LeakyRelu_l100_43_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_160) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43));
          end else begin
            if(when_LeakyRelu_l133_160) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_1));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_161) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_2));
          end else begin
            if(when_LeakyRelu_l133_161) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_3));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_162) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_4));
          end else begin
            if(when_LeakyRelu_l133_162) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_5));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_163) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_6));
          end else begin
            if(when_LeakyRelu_l133_163) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_7));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_164) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_8));
          end else begin
            if(when_LeakyRelu_l133_164) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_9));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_165) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_10));
          end else begin
            if(when_LeakyRelu_l133_165) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_11));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_166) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_12));
          end else begin
            if(when_LeakyRelu_l133_166) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_13));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_167) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_14));
          end else begin
            if(when_LeakyRelu_l133_167) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_15));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_168) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_16));
          end else begin
            if(when_LeakyRelu_l133_168) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_17));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_169) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_18));
          end else begin
            if(when_LeakyRelu_l133_169) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_19));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_170) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_20));
          end else begin
            if(when_LeakyRelu_l133_170) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_21));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_171) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_22));
          end else begin
            if(when_LeakyRelu_l133_171) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_23));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_172) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_24));
          end else begin
            if(when_LeakyRelu_l133_172) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_25));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_173) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_26));
          end else begin
            if(when_LeakyRelu_l133_173) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_27));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_174) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_28));
          end else begin
            if(when_LeakyRelu_l133_174) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_29));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_175) begin
            _zz_A_43 <= ($signed(_zz_A_40) + $signed(_zz__zz_A_43_30));
          end else begin
            if(when_LeakyRelu_l133_175) begin
              _zz_A_43 <= ($signed(_zz_A_40) - $signed(_zz__zz_A_43_31));
            end else begin
              _zz_A_43 <= _zz_A_40;
            end
          end
        end
        default : begin
          _zz_A_43 <= _zz_A_40;
        end
      endcase
    end else begin
      _zz_A_43 <= _zz_A_40;
    end
    if(when_LeakyRelu_l155_10) begin
      _zz_dataOut_10 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_10) begin
        _zz_dataOut_10 <= 8'hff;
      end else begin
        _zz_dataOut_10 <= _zz__zz_dataOut_10[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_45 <= _zz_when_LeakyRelu_l100_44;
    _zz_when_LeakyRelu_l100_46 <= _zz_when_LeakyRelu_l100_45;
    _zz_when_LeakyRelu_l100_47 <= _zz_when_LeakyRelu_l100_46;
    if(when_LeakyRelu_l100_11) begin
      if(when_LeakyRelu_l101_11) begin
        _zz_A_44 <= {{1{_zz_A_46[14]}}, _zz_A_46};
      end else begin
        if(when_LeakyRelu_l103_11) begin
          if(when_LeakyRelu_l104_11) begin
            _zz_A_44 <= {{1{_zz_A_45[14]}}, _zz_A_45};
          end else begin
            _zz_A_44 <= {{1{_zz_A_46[14]}}, _zz_A_46};
          end
        end else begin
          if(when_LeakyRelu_l110_11) begin
            _zz_A_44 <= {{1{_zz_A_45[14]}}, _zz_A_45};
          end else begin
            _zz_A_44 <= {{1{_zz_A_46[14]}}, _zz_A_46};
          end
        end
      end
    end else begin
      _zz_A_44 <= _zz_when_LeakyRelu_l100_47;
    end
    _zz_when_LeakyRelu_l100_47_regNext <= _zz_when_LeakyRelu_l100_47;
    if(when_LeakyRelu_l127_11) begin
      case(_zz_when_LeakyRelu_l100_47_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_176) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47));
          end else begin
            if(when_LeakyRelu_l133_176) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_1));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_177) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_2));
          end else begin
            if(when_LeakyRelu_l133_177) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_3));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_178) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_4));
          end else begin
            if(when_LeakyRelu_l133_178) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_5));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_179) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_6));
          end else begin
            if(when_LeakyRelu_l133_179) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_7));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_180) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_8));
          end else begin
            if(when_LeakyRelu_l133_180) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_9));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_181) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_10));
          end else begin
            if(when_LeakyRelu_l133_181) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_11));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_182) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_12));
          end else begin
            if(when_LeakyRelu_l133_182) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_13));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_183) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_14));
          end else begin
            if(when_LeakyRelu_l133_183) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_15));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_184) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_16));
          end else begin
            if(when_LeakyRelu_l133_184) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_17));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_185) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_18));
          end else begin
            if(when_LeakyRelu_l133_185) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_19));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_186) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_20));
          end else begin
            if(when_LeakyRelu_l133_186) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_21));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_187) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_22));
          end else begin
            if(when_LeakyRelu_l133_187) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_23));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_188) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_24));
          end else begin
            if(when_LeakyRelu_l133_188) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_25));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_189) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_26));
          end else begin
            if(when_LeakyRelu_l133_189) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_27));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_190) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_28));
          end else begin
            if(when_LeakyRelu_l133_190) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_29));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_191) begin
            _zz_A_47 <= ($signed(_zz_A_44) + $signed(_zz__zz_A_47_30));
          end else begin
            if(when_LeakyRelu_l133_191) begin
              _zz_A_47 <= ($signed(_zz_A_44) - $signed(_zz__zz_A_47_31));
            end else begin
              _zz_A_47 <= _zz_A_44;
            end
          end
        end
        default : begin
          _zz_A_47 <= _zz_A_44;
        end
      endcase
    end else begin
      _zz_A_47 <= _zz_A_44;
    end
    if(when_LeakyRelu_l155_11) begin
      _zz_dataOut_11 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_11) begin
        _zz_dataOut_11 <= 8'hff;
      end else begin
        _zz_dataOut_11 <= _zz__zz_dataOut_11[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_49 <= _zz_when_LeakyRelu_l100_48;
    _zz_when_LeakyRelu_l100_50 <= _zz_when_LeakyRelu_l100_49;
    _zz_when_LeakyRelu_l100_51 <= _zz_when_LeakyRelu_l100_50;
    if(when_LeakyRelu_l100_12) begin
      if(when_LeakyRelu_l101_12) begin
        _zz_A_48 <= {{1{_zz_A_50[14]}}, _zz_A_50};
      end else begin
        if(when_LeakyRelu_l103_12) begin
          if(when_LeakyRelu_l104_12) begin
            _zz_A_48 <= {{1{_zz_A_49[14]}}, _zz_A_49};
          end else begin
            _zz_A_48 <= {{1{_zz_A_50[14]}}, _zz_A_50};
          end
        end else begin
          if(when_LeakyRelu_l110_12) begin
            _zz_A_48 <= {{1{_zz_A_49[14]}}, _zz_A_49};
          end else begin
            _zz_A_48 <= {{1{_zz_A_50[14]}}, _zz_A_50};
          end
        end
      end
    end else begin
      _zz_A_48 <= _zz_when_LeakyRelu_l100_51;
    end
    _zz_when_LeakyRelu_l100_51_regNext <= _zz_when_LeakyRelu_l100_51;
    if(when_LeakyRelu_l127_12) begin
      case(_zz_when_LeakyRelu_l100_51_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_192) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51));
          end else begin
            if(when_LeakyRelu_l133_192) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_1));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_193) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_2));
          end else begin
            if(when_LeakyRelu_l133_193) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_3));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_194) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_4));
          end else begin
            if(when_LeakyRelu_l133_194) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_5));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_195) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_6));
          end else begin
            if(when_LeakyRelu_l133_195) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_7));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_196) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_8));
          end else begin
            if(when_LeakyRelu_l133_196) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_9));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_197) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_10));
          end else begin
            if(when_LeakyRelu_l133_197) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_11));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_198) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_12));
          end else begin
            if(when_LeakyRelu_l133_198) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_13));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_199) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_14));
          end else begin
            if(when_LeakyRelu_l133_199) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_15));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_200) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_16));
          end else begin
            if(when_LeakyRelu_l133_200) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_17));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_201) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_18));
          end else begin
            if(when_LeakyRelu_l133_201) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_19));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_202) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_20));
          end else begin
            if(when_LeakyRelu_l133_202) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_21));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_203) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_22));
          end else begin
            if(when_LeakyRelu_l133_203) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_23));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_204) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_24));
          end else begin
            if(when_LeakyRelu_l133_204) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_25));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_205) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_26));
          end else begin
            if(when_LeakyRelu_l133_205) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_27));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_206) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_28));
          end else begin
            if(when_LeakyRelu_l133_206) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_29));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_207) begin
            _zz_A_51 <= ($signed(_zz_A_48) + $signed(_zz__zz_A_51_30));
          end else begin
            if(when_LeakyRelu_l133_207) begin
              _zz_A_51 <= ($signed(_zz_A_48) - $signed(_zz__zz_A_51_31));
            end else begin
              _zz_A_51 <= _zz_A_48;
            end
          end
        end
        default : begin
          _zz_A_51 <= _zz_A_48;
        end
      endcase
    end else begin
      _zz_A_51 <= _zz_A_48;
    end
    if(when_LeakyRelu_l155_12) begin
      _zz_dataOut_12 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_12) begin
        _zz_dataOut_12 <= 8'hff;
      end else begin
        _zz_dataOut_12 <= _zz__zz_dataOut_12[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_53 <= _zz_when_LeakyRelu_l100_52;
    _zz_when_LeakyRelu_l100_54 <= _zz_when_LeakyRelu_l100_53;
    _zz_when_LeakyRelu_l100_55 <= _zz_when_LeakyRelu_l100_54;
    if(when_LeakyRelu_l100_13) begin
      if(when_LeakyRelu_l101_13) begin
        _zz_A_52 <= {{1{_zz_A_54[14]}}, _zz_A_54};
      end else begin
        if(when_LeakyRelu_l103_13) begin
          if(when_LeakyRelu_l104_13) begin
            _zz_A_52 <= {{1{_zz_A_53[14]}}, _zz_A_53};
          end else begin
            _zz_A_52 <= {{1{_zz_A_54[14]}}, _zz_A_54};
          end
        end else begin
          if(when_LeakyRelu_l110_13) begin
            _zz_A_52 <= {{1{_zz_A_53[14]}}, _zz_A_53};
          end else begin
            _zz_A_52 <= {{1{_zz_A_54[14]}}, _zz_A_54};
          end
        end
      end
    end else begin
      _zz_A_52 <= _zz_when_LeakyRelu_l100_55;
    end
    _zz_when_LeakyRelu_l100_55_regNext <= _zz_when_LeakyRelu_l100_55;
    if(when_LeakyRelu_l127_13) begin
      case(_zz_when_LeakyRelu_l100_55_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_208) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55));
          end else begin
            if(when_LeakyRelu_l133_208) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_1));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_209) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_2));
          end else begin
            if(when_LeakyRelu_l133_209) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_3));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_210) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_4));
          end else begin
            if(when_LeakyRelu_l133_210) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_5));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_211) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_6));
          end else begin
            if(when_LeakyRelu_l133_211) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_7));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_212) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_8));
          end else begin
            if(when_LeakyRelu_l133_212) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_9));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_213) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_10));
          end else begin
            if(when_LeakyRelu_l133_213) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_11));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_214) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_12));
          end else begin
            if(when_LeakyRelu_l133_214) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_13));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_215) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_14));
          end else begin
            if(when_LeakyRelu_l133_215) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_15));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_216) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_16));
          end else begin
            if(when_LeakyRelu_l133_216) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_17));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_217) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_18));
          end else begin
            if(when_LeakyRelu_l133_217) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_19));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_218) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_20));
          end else begin
            if(when_LeakyRelu_l133_218) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_21));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_219) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_22));
          end else begin
            if(when_LeakyRelu_l133_219) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_23));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_220) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_24));
          end else begin
            if(when_LeakyRelu_l133_220) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_25));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_221) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_26));
          end else begin
            if(when_LeakyRelu_l133_221) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_27));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_222) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_28));
          end else begin
            if(when_LeakyRelu_l133_222) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_29));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_223) begin
            _zz_A_55 <= ($signed(_zz_A_52) + $signed(_zz__zz_A_55_30));
          end else begin
            if(when_LeakyRelu_l133_223) begin
              _zz_A_55 <= ($signed(_zz_A_52) - $signed(_zz__zz_A_55_31));
            end else begin
              _zz_A_55 <= _zz_A_52;
            end
          end
        end
        default : begin
          _zz_A_55 <= _zz_A_52;
        end
      endcase
    end else begin
      _zz_A_55 <= _zz_A_52;
    end
    if(when_LeakyRelu_l155_13) begin
      _zz_dataOut_13 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_13) begin
        _zz_dataOut_13 <= 8'hff;
      end else begin
        _zz_dataOut_13 <= _zz__zz_dataOut_13[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_57 <= _zz_when_LeakyRelu_l100_56;
    _zz_when_LeakyRelu_l100_58 <= _zz_when_LeakyRelu_l100_57;
    _zz_when_LeakyRelu_l100_59 <= _zz_when_LeakyRelu_l100_58;
    if(when_LeakyRelu_l100_14) begin
      if(when_LeakyRelu_l101_14) begin
        _zz_A_56 <= {{1{_zz_A_58[14]}}, _zz_A_58};
      end else begin
        if(when_LeakyRelu_l103_14) begin
          if(when_LeakyRelu_l104_14) begin
            _zz_A_56 <= {{1{_zz_A_57[14]}}, _zz_A_57};
          end else begin
            _zz_A_56 <= {{1{_zz_A_58[14]}}, _zz_A_58};
          end
        end else begin
          if(when_LeakyRelu_l110_14) begin
            _zz_A_56 <= {{1{_zz_A_57[14]}}, _zz_A_57};
          end else begin
            _zz_A_56 <= {{1{_zz_A_58[14]}}, _zz_A_58};
          end
        end
      end
    end else begin
      _zz_A_56 <= _zz_when_LeakyRelu_l100_59;
    end
    _zz_when_LeakyRelu_l100_59_regNext <= _zz_when_LeakyRelu_l100_59;
    if(when_LeakyRelu_l127_14) begin
      case(_zz_when_LeakyRelu_l100_59_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_224) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59));
          end else begin
            if(when_LeakyRelu_l133_224) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_1));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_225) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_2));
          end else begin
            if(when_LeakyRelu_l133_225) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_3));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_226) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_4));
          end else begin
            if(when_LeakyRelu_l133_226) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_5));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_227) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_6));
          end else begin
            if(when_LeakyRelu_l133_227) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_7));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_228) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_8));
          end else begin
            if(when_LeakyRelu_l133_228) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_9));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_229) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_10));
          end else begin
            if(when_LeakyRelu_l133_229) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_11));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_230) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_12));
          end else begin
            if(when_LeakyRelu_l133_230) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_13));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_231) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_14));
          end else begin
            if(when_LeakyRelu_l133_231) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_15));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_232) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_16));
          end else begin
            if(when_LeakyRelu_l133_232) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_17));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_233) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_18));
          end else begin
            if(when_LeakyRelu_l133_233) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_19));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_234) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_20));
          end else begin
            if(when_LeakyRelu_l133_234) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_21));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_235) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_22));
          end else begin
            if(when_LeakyRelu_l133_235) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_23));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_236) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_24));
          end else begin
            if(when_LeakyRelu_l133_236) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_25));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_237) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_26));
          end else begin
            if(when_LeakyRelu_l133_237) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_27));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_238) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_28));
          end else begin
            if(when_LeakyRelu_l133_238) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_29));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_239) begin
            _zz_A_59 <= ($signed(_zz_A_56) + $signed(_zz__zz_A_59_30));
          end else begin
            if(when_LeakyRelu_l133_239) begin
              _zz_A_59 <= ($signed(_zz_A_56) - $signed(_zz__zz_A_59_31));
            end else begin
              _zz_A_59 <= _zz_A_56;
            end
          end
        end
        default : begin
          _zz_A_59 <= _zz_A_56;
        end
      endcase
    end else begin
      _zz_A_59 <= _zz_A_56;
    end
    if(when_LeakyRelu_l155_14) begin
      _zz_dataOut_14 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_14) begin
        _zz_dataOut_14 <= 8'hff;
      end else begin
        _zz_dataOut_14 <= _zz__zz_dataOut_14[7:0];
      end
    end
    _zz_when_LeakyRelu_l100_61 <= _zz_when_LeakyRelu_l100_60;
    _zz_when_LeakyRelu_l100_62 <= _zz_when_LeakyRelu_l100_61;
    _zz_when_LeakyRelu_l100_63 <= _zz_when_LeakyRelu_l100_62;
    if(when_LeakyRelu_l100_15) begin
      if(when_LeakyRelu_l101_15) begin
        _zz_A_60 <= {{1{_zz_A_62[14]}}, _zz_A_62};
      end else begin
        if(when_LeakyRelu_l103_15) begin
          if(when_LeakyRelu_l104_15) begin
            _zz_A_60 <= {{1{_zz_A_61[14]}}, _zz_A_61};
          end else begin
            _zz_A_60 <= {{1{_zz_A_62[14]}}, _zz_A_62};
          end
        end else begin
          if(when_LeakyRelu_l110_15) begin
            _zz_A_60 <= {{1{_zz_A_61[14]}}, _zz_A_61};
          end else begin
            _zz_A_60 <= {{1{_zz_A_62[14]}}, _zz_A_62};
          end
        end
      end
    end else begin
      _zz_A_60 <= _zz_when_LeakyRelu_l100_63;
    end
    _zz_when_LeakyRelu_l100_63_regNext <= _zz_when_LeakyRelu_l100_63;
    if(when_LeakyRelu_l127_15) begin
      case(_zz_when_LeakyRelu_l100_63_regNext)
        16'hfffb : begin
          if(when_LeakyRelu_l131_240) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63));
          end else begin
            if(when_LeakyRelu_l133_240) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_1));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hfff1 : begin
          if(when_LeakyRelu_l131_241) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_2));
          end else begin
            if(when_LeakyRelu_l133_241) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_3));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffe7 : begin
          if(when_LeakyRelu_l131_242) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_4));
          end else begin
            if(when_LeakyRelu_l133_242) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_5));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffdd : begin
          if(when_LeakyRelu_l131_243) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_6));
          end else begin
            if(when_LeakyRelu_l133_243) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_7));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffd3 : begin
          if(when_LeakyRelu_l131_244) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_8));
          end else begin
            if(when_LeakyRelu_l133_244) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_9));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffc9 : begin
          if(when_LeakyRelu_l131_245) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_10));
          end else begin
            if(when_LeakyRelu_l133_245) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_11));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffbf : begin
          if(when_LeakyRelu_l131_246) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_12));
          end else begin
            if(when_LeakyRelu_l133_246) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_13));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffb5 : begin
          if(when_LeakyRelu_l131_247) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_14));
          end else begin
            if(when_LeakyRelu_l133_247) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_15));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffab : begin
          if(when_LeakyRelu_l131_248) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_16));
          end else begin
            if(when_LeakyRelu_l133_248) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_17));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hffa1 : begin
          if(when_LeakyRelu_l131_249) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_18));
          end else begin
            if(when_LeakyRelu_l133_249) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_19));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff97 : begin
          if(when_LeakyRelu_l131_250) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_20));
          end else begin
            if(when_LeakyRelu_l133_250) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_21));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff8d : begin
          if(when_LeakyRelu_l131_251) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_22));
          end else begin
            if(when_LeakyRelu_l133_251) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_23));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff83 : begin
          if(when_LeakyRelu_l131_252) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_24));
          end else begin
            if(when_LeakyRelu_l133_252) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_25));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff79 : begin
          if(when_LeakyRelu_l131_253) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_26));
          end else begin
            if(when_LeakyRelu_l133_253) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_27));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff6f : begin
          if(when_LeakyRelu_l131_254) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_28));
          end else begin
            if(when_LeakyRelu_l133_254) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_29));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        16'hff65 : begin
          if(when_LeakyRelu_l131_255) begin
            _zz_A_63 <= ($signed(_zz_A_60) + $signed(_zz__zz_A_63_30));
          end else begin
            if(when_LeakyRelu_l133_255) begin
              _zz_A_63 <= ($signed(_zz_A_60) - $signed(_zz__zz_A_63_31));
            end else begin
              _zz_A_63 <= _zz_A_60;
            end
          end
        end
        default : begin
          _zz_A_63 <= _zz_A_60;
        end
      endcase
    end else begin
      _zz_A_63 <= _zz_A_60;
    end
    if(when_LeakyRelu_l155_15) begin
      _zz_dataOut_15 <= 8'h0;
    end else begin
      if(when_LeakyRelu_l157_15) begin
        _zz_dataOut_15 <= 8'hff;
      end else begin
        _zz_dataOut_15 <= _zz__zz_dataOut_15[7:0];
      end
    end
  end


endmodule

module Zero (
  input      [15:0]   dataIn_0,
  input      [15:0]   dataIn_1,
  input      [15:0]   dataIn_2,
  input      [15:0]   dataIn_3,
  input      [15:0]   dataIn_4,
  input      [15:0]   dataIn_5,
  input      [15:0]   dataIn_6,
  input      [15:0]   dataIn_7,
  input      [15:0]   dataIn_8,
  input      [15:0]   dataIn_9,
  input      [15:0]   dataIn_10,
  input      [15:0]   dataIn_11,
  input      [15:0]   dataIn_12,
  input      [15:0]   dataIn_13,
  input      [15:0]   dataIn_14,
  input      [15:0]   dataIn_15,
  input      [7:0]    quan_1,
  output     [7:0]    dataOut_0,
  output     [7:0]    dataOut_1,
  output     [7:0]    dataOut_2,
  output     [7:0]    dataOut_3,
  output     [7:0]    dataOut_4,
  output     [7:0]    dataOut_5,
  output     [7:0]    dataOut_6,
  output     [7:0]    dataOut_7,
  output     [7:0]    dataOut_8,
  output     [7:0]    dataOut_9,
  output     [7:0]    dataOut_10,
  output     [7:0]    dataOut_11,
  output     [7:0]    dataOut_12,
  output     [7:0]    dataOut_13,
  output     [7:0]    dataOut_14,
  output     [7:0]    dataOut_15,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [15:0]   addZero_0_S;
  wire       [15:0]   addZero_1_S;
  wire       [15:0]   addZero_2_S;
  wire       [15:0]   addZero_3_S;
  wire       [15:0]   addZero_4_S;
  wire       [15:0]   addZero_5_S;
  wire       [15:0]   addZero_6_S;
  wire       [15:0]   addZero_7_S;
  wire       [15:0]   addZero_8_S;
  wire       [15:0]   addZero_9_S;
  wire       [15:0]   addZero_10_S;
  wire       [15:0]   addZero_11_S;
  wire       [15:0]   addZero_12_S;
  wire       [15:0]   addZero_13_S;
  wire       [15:0]   addZero_14_S;
  wire       [15:0]   addZero_15_S;
  wire       [15:0]   _zz_normalData_0;
  wire       [15:0]   _zz_when_Quan_l173;
  wire       [15:0]   _zz_normalData_1;
  wire       [15:0]   _zz_when_Quan_l173_1;
  wire       [15:0]   _zz_normalData_2;
  wire       [15:0]   _zz_when_Quan_l173_2;
  wire       [15:0]   _zz_normalData_3;
  wire       [15:0]   _zz_when_Quan_l173_3;
  wire       [15:0]   _zz_normalData_4;
  wire       [15:0]   _zz_when_Quan_l173_4;
  wire       [15:0]   _zz_normalData_5;
  wire       [15:0]   _zz_when_Quan_l173_5;
  wire       [15:0]   _zz_normalData_6;
  wire       [15:0]   _zz_when_Quan_l173_6;
  wire       [15:0]   _zz_normalData_7;
  wire       [15:0]   _zz_when_Quan_l173_7;
  wire       [15:0]   _zz_normalData_8;
  wire       [15:0]   _zz_when_Quan_l173_8;
  wire       [15:0]   _zz_normalData_9;
  wire       [15:0]   _zz_when_Quan_l173_9;
  wire       [15:0]   _zz_normalData_10;
  wire       [15:0]   _zz_when_Quan_l173_10;
  wire       [15:0]   _zz_normalData_11;
  wire       [15:0]   _zz_when_Quan_l173_11;
  wire       [15:0]   _zz_normalData_12;
  wire       [15:0]   _zz_when_Quan_l173_12;
  wire       [15:0]   _zz_normalData_13;
  wire       [15:0]   _zz_when_Quan_l173_13;
  wire       [15:0]   _zz_normalData_14;
  wire       [15:0]   _zz_when_Quan_l173_14;
  wire       [15:0]   _zz_normalData_15;
  wire       [15:0]   _zz_when_Quan_l173_15;
  wire       [15:0]   addZeroTemp_0;
  wire       [15:0]   addZeroTemp_1;
  wire       [15:0]   addZeroTemp_2;
  wire       [15:0]   addZeroTemp_3;
  wire       [15:0]   addZeroTemp_4;
  wire       [15:0]   addZeroTemp_5;
  wire       [15:0]   addZeroTemp_6;
  wire       [15:0]   addZeroTemp_7;
  wire       [15:0]   addZeroTemp_8;
  wire       [15:0]   addZeroTemp_9;
  wire       [15:0]   addZeroTemp_10;
  wire       [15:0]   addZeroTemp_11;
  wire       [15:0]   addZeroTemp_12;
  wire       [15:0]   addZeroTemp_13;
  wire       [15:0]   addZeroTemp_14;
  wire       [15:0]   addZeroTemp_15;
  reg        [7:0]    normalData_0;
  reg        [7:0]    normalData_1;
  reg        [7:0]    normalData_2;
  reg        [7:0]    normalData_3;
  reg        [7:0]    normalData_4;
  reg        [7:0]    normalData_5;
  reg        [7:0]    normalData_6;
  reg        [7:0]    normalData_7;
  reg        [7:0]    normalData_8;
  reg        [7:0]    normalData_9;
  reg        [7:0]    normalData_10;
  reg        [7:0]    normalData_11;
  reg        [7:0]    normalData_12;
  reg        [7:0]    normalData_13;
  reg        [7:0]    normalData_14;
  reg        [7:0]    normalData_15;
  wire                when_Quan_l171;
  wire                when_Quan_l173;
  wire                when_Quan_l171_1;
  wire                when_Quan_l173_1;
  wire                when_Quan_l171_2;
  wire                when_Quan_l173_2;
  wire                when_Quan_l171_3;
  wire                when_Quan_l173_3;
  wire                when_Quan_l171_4;
  wire                when_Quan_l173_4;
  wire                when_Quan_l171_5;
  wire                when_Quan_l173_5;
  wire                when_Quan_l171_6;
  wire                when_Quan_l173_6;
  wire                when_Quan_l171_7;
  wire                when_Quan_l173_7;
  wire                when_Quan_l171_8;
  wire                when_Quan_l173_8;
  wire                when_Quan_l171_9;
  wire                when_Quan_l173_9;
  wire                when_Quan_l171_10;
  wire                when_Quan_l173_10;
  wire                when_Quan_l171_11;
  wire                when_Quan_l173_11;
  wire                when_Quan_l171_12;
  wire                when_Quan_l173_12;
  wire                when_Quan_l171_13;
  wire                when_Quan_l173_13;
  wire                when_Quan_l171_14;
  wire                when_Quan_l173_14;
  wire                when_Quan_l171_15;
  wire                when_Quan_l173_15;

  assign _zz_normalData_0 = addZeroTemp_0;
  assign _zz_when_Quan_l173 = 16'h00ff;
  assign _zz_normalData_1 = addZeroTemp_1;
  assign _zz_when_Quan_l173_1 = 16'h00ff;
  assign _zz_normalData_2 = addZeroTemp_2;
  assign _zz_when_Quan_l173_2 = 16'h00ff;
  assign _zz_normalData_3 = addZeroTemp_3;
  assign _zz_when_Quan_l173_3 = 16'h00ff;
  assign _zz_normalData_4 = addZeroTemp_4;
  assign _zz_when_Quan_l173_4 = 16'h00ff;
  assign _zz_normalData_5 = addZeroTemp_5;
  assign _zz_when_Quan_l173_5 = 16'h00ff;
  assign _zz_normalData_6 = addZeroTemp_6;
  assign _zz_when_Quan_l173_6 = 16'h00ff;
  assign _zz_normalData_7 = addZeroTemp_7;
  assign _zz_when_Quan_l173_7 = 16'h00ff;
  assign _zz_normalData_8 = addZeroTemp_8;
  assign _zz_when_Quan_l173_8 = 16'h00ff;
  assign _zz_normalData_9 = addZeroTemp_9;
  assign _zz_when_Quan_l173_9 = 16'h00ff;
  assign _zz_normalData_10 = addZeroTemp_10;
  assign _zz_when_Quan_l173_10 = 16'h00ff;
  assign _zz_normalData_11 = addZeroTemp_11;
  assign _zz_when_Quan_l173_11 = 16'h00ff;
  assign _zz_normalData_12 = addZeroTemp_12;
  assign _zz_when_Quan_l173_12 = 16'h00ff;
  assign _zz_normalData_13 = addZeroTemp_13;
  assign _zz_when_Quan_l173_13 = 16'h00ff;
  assign _zz_normalData_14 = addZeroTemp_14;
  assign _zz_when_Quan_l173_14 = 16'h00ff;
  assign _zz_normalData_15 = addZeroTemp_15;
  assign _zz_when_Quan_l173_15 = 16'h00ff;
  AddZero addZero_0 (
    .A   (dataIn_0[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_0_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_1 (
    .A   (dataIn_1[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_1_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_2 (
    .A   (dataIn_2[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_2_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_3 (
    .A   (dataIn_3[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_3_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_4 (
    .A   (dataIn_4[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_4_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_5 (
    .A   (dataIn_5[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_5_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_6 (
    .A   (dataIn_6[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_6_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_7 (
    .A   (dataIn_7[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_7_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_8 (
    .A   (dataIn_8[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_8_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_9 (
    .A   (dataIn_9[15:0]   ), //i
    .B   (quan_1[7:0]      ), //i
    .S   (addZero_9_S[15:0]), //o
    .CLK (clk              )  //i
  );
  AddZero addZero_10 (
    .A   (dataIn_10[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_10_S[15:0]), //o
    .CLK (clk               )  //i
  );
  AddZero addZero_11 (
    .A   (dataIn_11[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_11_S[15:0]), //o
    .CLK (clk               )  //i
  );
  AddZero addZero_12 (
    .A   (dataIn_12[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_12_S[15:0]), //o
    .CLK (clk               )  //i
  );
  AddZero addZero_13 (
    .A   (dataIn_13[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_13_S[15:0]), //o
    .CLK (clk               )  //i
  );
  AddZero addZero_14 (
    .A   (dataIn_14[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_14_S[15:0]), //o
    .CLK (clk               )  //i
  );
  AddZero addZero_15 (
    .A   (dataIn_15[15:0]   ), //i
    .B   (quan_1[7:0]       ), //i
    .S   (addZero_15_S[15:0]), //o
    .CLK (clk               )  //i
  );
  assign addZeroTemp_0 = addZero_0_S;
  assign addZeroTemp_1 = addZero_1_S;
  assign addZeroTemp_2 = addZero_2_S;
  assign addZeroTemp_3 = addZero_3_S;
  assign addZeroTemp_4 = addZero_4_S;
  assign addZeroTemp_5 = addZero_5_S;
  assign addZeroTemp_6 = addZero_6_S;
  assign addZeroTemp_7 = addZero_7_S;
  assign addZeroTemp_8 = addZero_8_S;
  assign addZeroTemp_9 = addZero_9_S;
  assign addZeroTemp_10 = addZero_10_S;
  assign addZeroTemp_11 = addZero_11_S;
  assign addZeroTemp_12 = addZero_12_S;
  assign addZeroTemp_13 = addZero_13_S;
  assign addZeroTemp_14 = addZero_14_S;
  assign addZeroTemp_15 = addZero_15_S;
  assign dataOut_0 = normalData_0;
  assign dataOut_1 = normalData_1;
  assign dataOut_2 = normalData_2;
  assign dataOut_3 = normalData_3;
  assign dataOut_4 = normalData_4;
  assign dataOut_5 = normalData_5;
  assign dataOut_6 = normalData_6;
  assign dataOut_7 = normalData_7;
  assign dataOut_8 = normalData_8;
  assign dataOut_9 = normalData_9;
  assign dataOut_10 = normalData_10;
  assign dataOut_11 = normalData_11;
  assign dataOut_12 = normalData_12;
  assign dataOut_13 = normalData_13;
  assign dataOut_14 = normalData_14;
  assign dataOut_15 = normalData_15;
  assign when_Quan_l171 = addZeroTemp_0[15];
  assign when_Quan_l173 = ($signed(_zz_when_Quan_l173) < $signed(addZeroTemp_0));
  assign when_Quan_l171_1 = addZeroTemp_1[15];
  assign when_Quan_l173_1 = ($signed(_zz_when_Quan_l173_1) < $signed(addZeroTemp_1));
  assign when_Quan_l171_2 = addZeroTemp_2[15];
  assign when_Quan_l173_2 = ($signed(_zz_when_Quan_l173_2) < $signed(addZeroTemp_2));
  assign when_Quan_l171_3 = addZeroTemp_3[15];
  assign when_Quan_l173_3 = ($signed(_zz_when_Quan_l173_3) < $signed(addZeroTemp_3));
  assign when_Quan_l171_4 = addZeroTemp_4[15];
  assign when_Quan_l173_4 = ($signed(_zz_when_Quan_l173_4) < $signed(addZeroTemp_4));
  assign when_Quan_l171_5 = addZeroTemp_5[15];
  assign when_Quan_l173_5 = ($signed(_zz_when_Quan_l173_5) < $signed(addZeroTemp_5));
  assign when_Quan_l171_6 = addZeroTemp_6[15];
  assign when_Quan_l173_6 = ($signed(_zz_when_Quan_l173_6) < $signed(addZeroTemp_6));
  assign when_Quan_l171_7 = addZeroTemp_7[15];
  assign when_Quan_l173_7 = ($signed(_zz_when_Quan_l173_7) < $signed(addZeroTemp_7));
  assign when_Quan_l171_8 = addZeroTemp_8[15];
  assign when_Quan_l173_8 = ($signed(_zz_when_Quan_l173_8) < $signed(addZeroTemp_8));
  assign when_Quan_l171_9 = addZeroTemp_9[15];
  assign when_Quan_l173_9 = ($signed(_zz_when_Quan_l173_9) < $signed(addZeroTemp_9));
  assign when_Quan_l171_10 = addZeroTemp_10[15];
  assign when_Quan_l173_10 = ($signed(_zz_when_Quan_l173_10) < $signed(addZeroTemp_10));
  assign when_Quan_l171_11 = addZeroTemp_11[15];
  assign when_Quan_l173_11 = ($signed(_zz_when_Quan_l173_11) < $signed(addZeroTemp_11));
  assign when_Quan_l171_12 = addZeroTemp_12[15];
  assign when_Quan_l173_12 = ($signed(_zz_when_Quan_l173_12) < $signed(addZeroTemp_12));
  assign when_Quan_l171_13 = addZeroTemp_13[15];
  assign when_Quan_l173_13 = ($signed(_zz_when_Quan_l173_13) < $signed(addZeroTemp_13));
  assign when_Quan_l171_14 = addZeroTemp_14[15];
  assign when_Quan_l173_14 = ($signed(_zz_when_Quan_l173_14) < $signed(addZeroTemp_14));
  assign when_Quan_l171_15 = addZeroTemp_15[15];
  assign when_Quan_l173_15 = ($signed(_zz_when_Quan_l173_15) < $signed(addZeroTemp_15));
  always @(posedge clk) begin
    if(when_Quan_l171) begin
      normalData_0 <= 8'h0;
    end else begin
      if(when_Quan_l173) begin
        normalData_0 <= 8'hff;
      end else begin
        normalData_0 <= _zz_normalData_0[7:0];
      end
    end
    if(when_Quan_l171_1) begin
      normalData_1 <= 8'h0;
    end else begin
      if(when_Quan_l173_1) begin
        normalData_1 <= 8'hff;
      end else begin
        normalData_1 <= _zz_normalData_1[7:0];
      end
    end
    if(when_Quan_l171_2) begin
      normalData_2 <= 8'h0;
    end else begin
      if(when_Quan_l173_2) begin
        normalData_2 <= 8'hff;
      end else begin
        normalData_2 <= _zz_normalData_2[7:0];
      end
    end
    if(when_Quan_l171_3) begin
      normalData_3 <= 8'h0;
    end else begin
      if(when_Quan_l173_3) begin
        normalData_3 <= 8'hff;
      end else begin
        normalData_3 <= _zz_normalData_3[7:0];
      end
    end
    if(when_Quan_l171_4) begin
      normalData_4 <= 8'h0;
    end else begin
      if(when_Quan_l173_4) begin
        normalData_4 <= 8'hff;
      end else begin
        normalData_4 <= _zz_normalData_4[7:0];
      end
    end
    if(when_Quan_l171_5) begin
      normalData_5 <= 8'h0;
    end else begin
      if(when_Quan_l173_5) begin
        normalData_5 <= 8'hff;
      end else begin
        normalData_5 <= _zz_normalData_5[7:0];
      end
    end
    if(when_Quan_l171_6) begin
      normalData_6 <= 8'h0;
    end else begin
      if(when_Quan_l173_6) begin
        normalData_6 <= 8'hff;
      end else begin
        normalData_6 <= _zz_normalData_6[7:0];
      end
    end
    if(when_Quan_l171_7) begin
      normalData_7 <= 8'h0;
    end else begin
      if(when_Quan_l173_7) begin
        normalData_7 <= 8'hff;
      end else begin
        normalData_7 <= _zz_normalData_7[7:0];
      end
    end
    if(when_Quan_l171_8) begin
      normalData_8 <= 8'h0;
    end else begin
      if(when_Quan_l173_8) begin
        normalData_8 <= 8'hff;
      end else begin
        normalData_8 <= _zz_normalData_8[7:0];
      end
    end
    if(when_Quan_l171_9) begin
      normalData_9 <= 8'h0;
    end else begin
      if(when_Quan_l173_9) begin
        normalData_9 <= 8'hff;
      end else begin
        normalData_9 <= _zz_normalData_9[7:0];
      end
    end
    if(when_Quan_l171_10) begin
      normalData_10 <= 8'h0;
    end else begin
      if(when_Quan_l173_10) begin
        normalData_10 <= 8'hff;
      end else begin
        normalData_10 <= _zz_normalData_10[7:0];
      end
    end
    if(when_Quan_l171_11) begin
      normalData_11 <= 8'h0;
    end else begin
      if(when_Quan_l173_11) begin
        normalData_11 <= 8'hff;
      end else begin
        normalData_11 <= _zz_normalData_11[7:0];
      end
    end
    if(when_Quan_l171_12) begin
      normalData_12 <= 8'h0;
    end else begin
      if(when_Quan_l173_12) begin
        normalData_12 <= 8'hff;
      end else begin
        normalData_12 <= _zz_normalData_12[7:0];
      end
    end
    if(when_Quan_l171_13) begin
      normalData_13 <= 8'h0;
    end else begin
      if(when_Quan_l173_13) begin
        normalData_13 <= 8'hff;
      end else begin
        normalData_13 <= _zz_normalData_13[7:0];
      end
    end
    if(when_Quan_l171_14) begin
      normalData_14 <= 8'h0;
    end else begin
      if(when_Quan_l173_14) begin
        normalData_14 <= 8'hff;
      end else begin
        normalData_14 <= _zz_normalData_14[7:0];
      end
    end
    if(when_Quan_l171_15) begin
      normalData_15 <= 8'h0;
    end else begin
      if(when_Quan_l173_15) begin
        normalData_15 <= 8'hff;
      end else begin
        normalData_15 <= _zz_normalData_15[7:0];
      end
    end
  end


endmodule

module Shift (
  input      [31:0]   shift_dataIn_0,
  input      [31:0]   shift_dataIn_1,
  input      [31:0]   shift_dataIn_2,
  input      [31:0]   shift_dataIn_3,
  input      [31:0]   shift_dataIn_4,
  input      [31:0]   shift_dataIn_5,
  input      [31:0]   shift_dataIn_6,
  input      [31:0]   shift_dataIn_7,
  input      [31:0]   shift_dataIn_8,
  input      [31:0]   shift_dataIn_9,
  input      [31:0]   shift_dataIn_10,
  input      [31:0]   shift_dataIn_11,
  input      [31:0]   shift_dataIn_12,
  input      [31:0]   shift_dataIn_13,
  input      [31:0]   shift_dataIn_14,
  input      [31:0]   shift_dataIn_15,
  input      [31:0]   shift_quan_0,
  input      [31:0]   shift_quan_1,
  input      [31:0]   shift_quan_2,
  input      [31:0]   shift_quan_3,
  input      [31:0]   shift_quan_4,
  input      [31:0]   shift_quan_5,
  input      [31:0]   shift_quan_6,
  input      [31:0]   shift_quan_7,
  input      [31:0]   shift_quan_8,
  input      [31:0]   shift_quan_9,
  input      [31:0]   shift_quan_10,
  input      [31:0]   shift_quan_11,
  input      [31:0]   shift_quan_12,
  input      [31:0]   shift_quan_13,
  input      [31:0]   shift_quan_14,
  input      [31:0]   shift_quan_15,
  output     [15:0]   shift_dataOut_0,
  output     [15:0]   shift_dataOut_1,
  output     [15:0]   shift_dataOut_2,
  output     [15:0]   shift_dataOut_3,
  output     [15:0]   shift_dataOut_4,
  output     [15:0]   shift_dataOut_5,
  output     [15:0]   shift_dataOut_6,
  output     [15:0]   shift_dataOut_7,
  output     [15:0]   shift_dataOut_8,
  output     [15:0]   shift_dataOut_9,
  output     [15:0]   shift_dataOut_10,
  output     [15:0]   shift_dataOut_11,
  output     [15:0]   shift_dataOut_12,
  output     [15:0]   shift_dataOut_13,
  output     [15:0]   shift_dataOut_14,
  output     [15:0]   shift_dataOut_15,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [15:0]   _zz__zz_shift_dataOut_0_1;
  wire       [0:0]    _zz__zz_shift_dataOut_0_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_0_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_0_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_0_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_0_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_1_1;
  wire       [0:0]    _zz__zz_shift_dataOut_1_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_1_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_1_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_1_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_1_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_2_1;
  wire       [0:0]    _zz__zz_shift_dataOut_2_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_2_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_2_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_2_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_2_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_3_1;
  wire       [0:0]    _zz__zz_shift_dataOut_3_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_3_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_3_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_3_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_3_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_4_1;
  wire       [0:0]    _zz__zz_shift_dataOut_4_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_4_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_4_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_4_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_4_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_5_1;
  wire       [0:0]    _zz__zz_shift_dataOut_5_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_5_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_5_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_5_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_5_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_6_1;
  wire       [0:0]    _zz__zz_shift_dataOut_6_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_6_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_6_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_6_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_6_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_7_1;
  wire       [0:0]    _zz__zz_shift_dataOut_7_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_7_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_7_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_7_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_7_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_8_1;
  wire       [0:0]    _zz__zz_shift_dataOut_8_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_8_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_8_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_8_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_8_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_9_1;
  wire       [0:0]    _zz__zz_shift_dataOut_9_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_9_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_9_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_9_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_9_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_10_1;
  wire       [0:0]    _zz__zz_shift_dataOut_10_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_10_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_10_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_10_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_10_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_11_1;
  wire       [0:0]    _zz__zz_shift_dataOut_11_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_11_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_11_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_11_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_11_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_12_1;
  wire       [0:0]    _zz__zz_shift_dataOut_12_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_12_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_12_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_12_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_12_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_13_1;
  wire       [0:0]    _zz__zz_shift_dataOut_13_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_13_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_13_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_13_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_13_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_14_1;
  wire       [0:0]    _zz__zz_shift_dataOut_14_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_14_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_14_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_14_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_14_1_5;
  wire       [15:0]   _zz__zz_shift_dataOut_15_1;
  wire       [0:0]    _zz__zz_shift_dataOut_15_1_1;
  wire       [14:0]   _zz__zz_shift_dataOut_15_1_2;
  wire       [15:0]   _zz__zz_shift_dataOut_15_1_3;
  wire       [0:0]    _zz__zz_shift_dataOut_15_1_4;
  wire       [14:0]   _zz__zz_shift_dataOut_15_1_5;
  wire       [31:0]   _zz_shift_dataOut_0;
  reg        [15:0]   _zz_shift_dataOut_0_1;
  wire                when_Quan_l130;
  wire       [31:0]   _zz_shift_dataOut_1;
  reg        [15:0]   _zz_shift_dataOut_1_1;
  wire                when_Quan_l130_1;
  wire       [31:0]   _zz_shift_dataOut_2;
  reg        [15:0]   _zz_shift_dataOut_2_1;
  wire                when_Quan_l130_2;
  wire       [31:0]   _zz_shift_dataOut_3;
  reg        [15:0]   _zz_shift_dataOut_3_1;
  wire                when_Quan_l130_3;
  wire       [31:0]   _zz_shift_dataOut_4;
  reg        [15:0]   _zz_shift_dataOut_4_1;
  wire                when_Quan_l130_4;
  wire       [31:0]   _zz_shift_dataOut_5;
  reg        [15:0]   _zz_shift_dataOut_5_1;
  wire                when_Quan_l130_5;
  wire       [31:0]   _zz_shift_dataOut_6;
  reg        [15:0]   _zz_shift_dataOut_6_1;
  wire                when_Quan_l130_6;
  wire       [31:0]   _zz_shift_dataOut_7;
  reg        [15:0]   _zz_shift_dataOut_7_1;
  wire                when_Quan_l130_7;
  wire       [31:0]   _zz_shift_dataOut_8;
  reg        [15:0]   _zz_shift_dataOut_8_1;
  wire                when_Quan_l130_8;
  wire       [31:0]   _zz_shift_dataOut_9;
  reg        [15:0]   _zz_shift_dataOut_9_1;
  wire                when_Quan_l130_9;
  wire       [31:0]   _zz_shift_dataOut_10;
  reg        [15:0]   _zz_shift_dataOut_10_1;
  wire                when_Quan_l130_10;
  wire       [31:0]   _zz_shift_dataOut_11;
  reg        [15:0]   _zz_shift_dataOut_11_1;
  wire                when_Quan_l130_11;
  wire       [31:0]   _zz_shift_dataOut_12;
  reg        [15:0]   _zz_shift_dataOut_12_1;
  wire                when_Quan_l130_12;
  wire       [31:0]   _zz_shift_dataOut_13;
  reg        [15:0]   _zz_shift_dataOut_13_1;
  wire                when_Quan_l130_13;
  wire       [31:0]   _zz_shift_dataOut_14;
  reg        [15:0]   _zz_shift_dataOut_14_1;
  wire                when_Quan_l130_14;
  wire       [31:0]   _zz_shift_dataOut_15;
  reg        [15:0]   _zz_shift_dataOut_15_1;
  wire                when_Quan_l130_15;

  assign _zz__zz_shift_dataOut_0_1 = {_zz__zz_shift_dataOut_0_1_1,_zz__zz_shift_dataOut_0_1_2};
  assign _zz__zz_shift_dataOut_0_1_1 = _zz_shift_dataOut_0[31];
  assign _zz__zz_shift_dataOut_0_1_2 = _zz_shift_dataOut_0[15 : 1];
  assign _zz__zz_shift_dataOut_0_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_0_1_4 = _zz_shift_dataOut_0[31];
  assign _zz__zz_shift_dataOut_0_1_5 = _zz_shift_dataOut_0[15 : 1];
  assign _zz__zz_shift_dataOut_1_1 = {_zz__zz_shift_dataOut_1_1_1,_zz__zz_shift_dataOut_1_1_2};
  assign _zz__zz_shift_dataOut_1_1_1 = _zz_shift_dataOut_1[31];
  assign _zz__zz_shift_dataOut_1_1_2 = _zz_shift_dataOut_1[15 : 1];
  assign _zz__zz_shift_dataOut_1_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_1_1_4 = _zz_shift_dataOut_1[31];
  assign _zz__zz_shift_dataOut_1_1_5 = _zz_shift_dataOut_1[15 : 1];
  assign _zz__zz_shift_dataOut_2_1 = {_zz__zz_shift_dataOut_2_1_1,_zz__zz_shift_dataOut_2_1_2};
  assign _zz__zz_shift_dataOut_2_1_1 = _zz_shift_dataOut_2[31];
  assign _zz__zz_shift_dataOut_2_1_2 = _zz_shift_dataOut_2[15 : 1];
  assign _zz__zz_shift_dataOut_2_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_2_1_4 = _zz_shift_dataOut_2[31];
  assign _zz__zz_shift_dataOut_2_1_5 = _zz_shift_dataOut_2[15 : 1];
  assign _zz__zz_shift_dataOut_3_1 = {_zz__zz_shift_dataOut_3_1_1,_zz__zz_shift_dataOut_3_1_2};
  assign _zz__zz_shift_dataOut_3_1_1 = _zz_shift_dataOut_3[31];
  assign _zz__zz_shift_dataOut_3_1_2 = _zz_shift_dataOut_3[15 : 1];
  assign _zz__zz_shift_dataOut_3_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_3_1_4 = _zz_shift_dataOut_3[31];
  assign _zz__zz_shift_dataOut_3_1_5 = _zz_shift_dataOut_3[15 : 1];
  assign _zz__zz_shift_dataOut_4_1 = {_zz__zz_shift_dataOut_4_1_1,_zz__zz_shift_dataOut_4_1_2};
  assign _zz__zz_shift_dataOut_4_1_1 = _zz_shift_dataOut_4[31];
  assign _zz__zz_shift_dataOut_4_1_2 = _zz_shift_dataOut_4[15 : 1];
  assign _zz__zz_shift_dataOut_4_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_4_1_4 = _zz_shift_dataOut_4[31];
  assign _zz__zz_shift_dataOut_4_1_5 = _zz_shift_dataOut_4[15 : 1];
  assign _zz__zz_shift_dataOut_5_1 = {_zz__zz_shift_dataOut_5_1_1,_zz__zz_shift_dataOut_5_1_2};
  assign _zz__zz_shift_dataOut_5_1_1 = _zz_shift_dataOut_5[31];
  assign _zz__zz_shift_dataOut_5_1_2 = _zz_shift_dataOut_5[15 : 1];
  assign _zz__zz_shift_dataOut_5_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_5_1_4 = _zz_shift_dataOut_5[31];
  assign _zz__zz_shift_dataOut_5_1_5 = _zz_shift_dataOut_5[15 : 1];
  assign _zz__zz_shift_dataOut_6_1 = {_zz__zz_shift_dataOut_6_1_1,_zz__zz_shift_dataOut_6_1_2};
  assign _zz__zz_shift_dataOut_6_1_1 = _zz_shift_dataOut_6[31];
  assign _zz__zz_shift_dataOut_6_1_2 = _zz_shift_dataOut_6[15 : 1];
  assign _zz__zz_shift_dataOut_6_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_6_1_4 = _zz_shift_dataOut_6[31];
  assign _zz__zz_shift_dataOut_6_1_5 = _zz_shift_dataOut_6[15 : 1];
  assign _zz__zz_shift_dataOut_7_1 = {_zz__zz_shift_dataOut_7_1_1,_zz__zz_shift_dataOut_7_1_2};
  assign _zz__zz_shift_dataOut_7_1_1 = _zz_shift_dataOut_7[31];
  assign _zz__zz_shift_dataOut_7_1_2 = _zz_shift_dataOut_7[15 : 1];
  assign _zz__zz_shift_dataOut_7_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_7_1_4 = _zz_shift_dataOut_7[31];
  assign _zz__zz_shift_dataOut_7_1_5 = _zz_shift_dataOut_7[15 : 1];
  assign _zz__zz_shift_dataOut_8_1 = {_zz__zz_shift_dataOut_8_1_1,_zz__zz_shift_dataOut_8_1_2};
  assign _zz__zz_shift_dataOut_8_1_1 = _zz_shift_dataOut_8[31];
  assign _zz__zz_shift_dataOut_8_1_2 = _zz_shift_dataOut_8[15 : 1];
  assign _zz__zz_shift_dataOut_8_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_8_1_4 = _zz_shift_dataOut_8[31];
  assign _zz__zz_shift_dataOut_8_1_5 = _zz_shift_dataOut_8[15 : 1];
  assign _zz__zz_shift_dataOut_9_1 = {_zz__zz_shift_dataOut_9_1_1,_zz__zz_shift_dataOut_9_1_2};
  assign _zz__zz_shift_dataOut_9_1_1 = _zz_shift_dataOut_9[31];
  assign _zz__zz_shift_dataOut_9_1_2 = _zz_shift_dataOut_9[15 : 1];
  assign _zz__zz_shift_dataOut_9_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_9_1_4 = _zz_shift_dataOut_9[31];
  assign _zz__zz_shift_dataOut_9_1_5 = _zz_shift_dataOut_9[15 : 1];
  assign _zz__zz_shift_dataOut_10_1 = {_zz__zz_shift_dataOut_10_1_1,_zz__zz_shift_dataOut_10_1_2};
  assign _zz__zz_shift_dataOut_10_1_1 = _zz_shift_dataOut_10[31];
  assign _zz__zz_shift_dataOut_10_1_2 = _zz_shift_dataOut_10[15 : 1];
  assign _zz__zz_shift_dataOut_10_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_10_1_4 = _zz_shift_dataOut_10[31];
  assign _zz__zz_shift_dataOut_10_1_5 = _zz_shift_dataOut_10[15 : 1];
  assign _zz__zz_shift_dataOut_11_1 = {_zz__zz_shift_dataOut_11_1_1,_zz__zz_shift_dataOut_11_1_2};
  assign _zz__zz_shift_dataOut_11_1_1 = _zz_shift_dataOut_11[31];
  assign _zz__zz_shift_dataOut_11_1_2 = _zz_shift_dataOut_11[15 : 1];
  assign _zz__zz_shift_dataOut_11_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_11_1_4 = _zz_shift_dataOut_11[31];
  assign _zz__zz_shift_dataOut_11_1_5 = _zz_shift_dataOut_11[15 : 1];
  assign _zz__zz_shift_dataOut_12_1 = {_zz__zz_shift_dataOut_12_1_1,_zz__zz_shift_dataOut_12_1_2};
  assign _zz__zz_shift_dataOut_12_1_1 = _zz_shift_dataOut_12[31];
  assign _zz__zz_shift_dataOut_12_1_2 = _zz_shift_dataOut_12[15 : 1];
  assign _zz__zz_shift_dataOut_12_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_12_1_4 = _zz_shift_dataOut_12[31];
  assign _zz__zz_shift_dataOut_12_1_5 = _zz_shift_dataOut_12[15 : 1];
  assign _zz__zz_shift_dataOut_13_1 = {_zz__zz_shift_dataOut_13_1_1,_zz__zz_shift_dataOut_13_1_2};
  assign _zz__zz_shift_dataOut_13_1_1 = _zz_shift_dataOut_13[31];
  assign _zz__zz_shift_dataOut_13_1_2 = _zz_shift_dataOut_13[15 : 1];
  assign _zz__zz_shift_dataOut_13_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_13_1_4 = _zz_shift_dataOut_13[31];
  assign _zz__zz_shift_dataOut_13_1_5 = _zz_shift_dataOut_13[15 : 1];
  assign _zz__zz_shift_dataOut_14_1 = {_zz__zz_shift_dataOut_14_1_1,_zz__zz_shift_dataOut_14_1_2};
  assign _zz__zz_shift_dataOut_14_1_1 = _zz_shift_dataOut_14[31];
  assign _zz__zz_shift_dataOut_14_1_2 = _zz_shift_dataOut_14[15 : 1];
  assign _zz__zz_shift_dataOut_14_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_14_1_4 = _zz_shift_dataOut_14[31];
  assign _zz__zz_shift_dataOut_14_1_5 = _zz_shift_dataOut_14[15 : 1];
  assign _zz__zz_shift_dataOut_15_1 = {_zz__zz_shift_dataOut_15_1_1,_zz__zz_shift_dataOut_15_1_2};
  assign _zz__zz_shift_dataOut_15_1_1 = _zz_shift_dataOut_15[31];
  assign _zz__zz_shift_dataOut_15_1_2 = _zz_shift_dataOut_15[15 : 1];
  assign _zz__zz_shift_dataOut_15_1_3 = 16'h0001;
  assign _zz__zz_shift_dataOut_15_1_4 = _zz_shift_dataOut_15[31];
  assign _zz__zz_shift_dataOut_15_1_5 = _zz_shift_dataOut_15[15 : 1];
  assign _zz_shift_dataOut_0 = ($signed(shift_dataIn_0) >>> shift_quan_0);
  assign when_Quan_l130 = _zz_shift_dataOut_0[0];
  assign shift_dataOut_0 = _zz_shift_dataOut_0_1;
  assign _zz_shift_dataOut_1 = ($signed(shift_dataIn_1) >>> shift_quan_1);
  assign when_Quan_l130_1 = _zz_shift_dataOut_1[0];
  assign shift_dataOut_1 = _zz_shift_dataOut_1_1;
  assign _zz_shift_dataOut_2 = ($signed(shift_dataIn_2) >>> shift_quan_2);
  assign when_Quan_l130_2 = _zz_shift_dataOut_2[0];
  assign shift_dataOut_2 = _zz_shift_dataOut_2_1;
  assign _zz_shift_dataOut_3 = ($signed(shift_dataIn_3) >>> shift_quan_3);
  assign when_Quan_l130_3 = _zz_shift_dataOut_3[0];
  assign shift_dataOut_3 = _zz_shift_dataOut_3_1;
  assign _zz_shift_dataOut_4 = ($signed(shift_dataIn_4) >>> shift_quan_4);
  assign when_Quan_l130_4 = _zz_shift_dataOut_4[0];
  assign shift_dataOut_4 = _zz_shift_dataOut_4_1;
  assign _zz_shift_dataOut_5 = ($signed(shift_dataIn_5) >>> shift_quan_5);
  assign when_Quan_l130_5 = _zz_shift_dataOut_5[0];
  assign shift_dataOut_5 = _zz_shift_dataOut_5_1;
  assign _zz_shift_dataOut_6 = ($signed(shift_dataIn_6) >>> shift_quan_6);
  assign when_Quan_l130_6 = _zz_shift_dataOut_6[0];
  assign shift_dataOut_6 = _zz_shift_dataOut_6_1;
  assign _zz_shift_dataOut_7 = ($signed(shift_dataIn_7) >>> shift_quan_7);
  assign when_Quan_l130_7 = _zz_shift_dataOut_7[0];
  assign shift_dataOut_7 = _zz_shift_dataOut_7_1;
  assign _zz_shift_dataOut_8 = ($signed(shift_dataIn_8) >>> shift_quan_8);
  assign when_Quan_l130_8 = _zz_shift_dataOut_8[0];
  assign shift_dataOut_8 = _zz_shift_dataOut_8_1;
  assign _zz_shift_dataOut_9 = ($signed(shift_dataIn_9) >>> shift_quan_9);
  assign when_Quan_l130_9 = _zz_shift_dataOut_9[0];
  assign shift_dataOut_9 = _zz_shift_dataOut_9_1;
  assign _zz_shift_dataOut_10 = ($signed(shift_dataIn_10) >>> shift_quan_10);
  assign when_Quan_l130_10 = _zz_shift_dataOut_10[0];
  assign shift_dataOut_10 = _zz_shift_dataOut_10_1;
  assign _zz_shift_dataOut_11 = ($signed(shift_dataIn_11) >>> shift_quan_11);
  assign when_Quan_l130_11 = _zz_shift_dataOut_11[0];
  assign shift_dataOut_11 = _zz_shift_dataOut_11_1;
  assign _zz_shift_dataOut_12 = ($signed(shift_dataIn_12) >>> shift_quan_12);
  assign when_Quan_l130_12 = _zz_shift_dataOut_12[0];
  assign shift_dataOut_12 = _zz_shift_dataOut_12_1;
  assign _zz_shift_dataOut_13 = ($signed(shift_dataIn_13) >>> shift_quan_13);
  assign when_Quan_l130_13 = _zz_shift_dataOut_13[0];
  assign shift_dataOut_13 = _zz_shift_dataOut_13_1;
  assign _zz_shift_dataOut_14 = ($signed(shift_dataIn_14) >>> shift_quan_14);
  assign when_Quan_l130_14 = _zz_shift_dataOut_14[0];
  assign shift_dataOut_14 = _zz_shift_dataOut_14_1;
  assign _zz_shift_dataOut_15 = ($signed(shift_dataIn_15) >>> shift_quan_15);
  assign when_Quan_l130_15 = _zz_shift_dataOut_15[0];
  assign shift_dataOut_15 = _zz_shift_dataOut_15_1;
  always @(posedge clk) begin
    if(when_Quan_l130) begin
      _zz_shift_dataOut_0_1 <= ($signed(_zz__zz_shift_dataOut_0_1) + $signed(_zz__zz_shift_dataOut_0_1_3));
    end else begin
      _zz_shift_dataOut_0_1 <= {_zz__zz_shift_dataOut_0_1_4,_zz__zz_shift_dataOut_0_1_5};
    end
    if(when_Quan_l130_1) begin
      _zz_shift_dataOut_1_1 <= ($signed(_zz__zz_shift_dataOut_1_1) + $signed(_zz__zz_shift_dataOut_1_1_3));
    end else begin
      _zz_shift_dataOut_1_1 <= {_zz__zz_shift_dataOut_1_1_4,_zz__zz_shift_dataOut_1_1_5};
    end
    if(when_Quan_l130_2) begin
      _zz_shift_dataOut_2_1 <= ($signed(_zz__zz_shift_dataOut_2_1) + $signed(_zz__zz_shift_dataOut_2_1_3));
    end else begin
      _zz_shift_dataOut_2_1 <= {_zz__zz_shift_dataOut_2_1_4,_zz__zz_shift_dataOut_2_1_5};
    end
    if(when_Quan_l130_3) begin
      _zz_shift_dataOut_3_1 <= ($signed(_zz__zz_shift_dataOut_3_1) + $signed(_zz__zz_shift_dataOut_3_1_3));
    end else begin
      _zz_shift_dataOut_3_1 <= {_zz__zz_shift_dataOut_3_1_4,_zz__zz_shift_dataOut_3_1_5};
    end
    if(when_Quan_l130_4) begin
      _zz_shift_dataOut_4_1 <= ($signed(_zz__zz_shift_dataOut_4_1) + $signed(_zz__zz_shift_dataOut_4_1_3));
    end else begin
      _zz_shift_dataOut_4_1 <= {_zz__zz_shift_dataOut_4_1_4,_zz__zz_shift_dataOut_4_1_5};
    end
    if(when_Quan_l130_5) begin
      _zz_shift_dataOut_5_1 <= ($signed(_zz__zz_shift_dataOut_5_1) + $signed(_zz__zz_shift_dataOut_5_1_3));
    end else begin
      _zz_shift_dataOut_5_1 <= {_zz__zz_shift_dataOut_5_1_4,_zz__zz_shift_dataOut_5_1_5};
    end
    if(when_Quan_l130_6) begin
      _zz_shift_dataOut_6_1 <= ($signed(_zz__zz_shift_dataOut_6_1) + $signed(_zz__zz_shift_dataOut_6_1_3));
    end else begin
      _zz_shift_dataOut_6_1 <= {_zz__zz_shift_dataOut_6_1_4,_zz__zz_shift_dataOut_6_1_5};
    end
    if(when_Quan_l130_7) begin
      _zz_shift_dataOut_7_1 <= ($signed(_zz__zz_shift_dataOut_7_1) + $signed(_zz__zz_shift_dataOut_7_1_3));
    end else begin
      _zz_shift_dataOut_7_1 <= {_zz__zz_shift_dataOut_7_1_4,_zz__zz_shift_dataOut_7_1_5};
    end
    if(when_Quan_l130_8) begin
      _zz_shift_dataOut_8_1 <= ($signed(_zz__zz_shift_dataOut_8_1) + $signed(_zz__zz_shift_dataOut_8_1_3));
    end else begin
      _zz_shift_dataOut_8_1 <= {_zz__zz_shift_dataOut_8_1_4,_zz__zz_shift_dataOut_8_1_5};
    end
    if(when_Quan_l130_9) begin
      _zz_shift_dataOut_9_1 <= ($signed(_zz__zz_shift_dataOut_9_1) + $signed(_zz__zz_shift_dataOut_9_1_3));
    end else begin
      _zz_shift_dataOut_9_1 <= {_zz__zz_shift_dataOut_9_1_4,_zz__zz_shift_dataOut_9_1_5};
    end
    if(when_Quan_l130_10) begin
      _zz_shift_dataOut_10_1 <= ($signed(_zz__zz_shift_dataOut_10_1) + $signed(_zz__zz_shift_dataOut_10_1_3));
    end else begin
      _zz_shift_dataOut_10_1 <= {_zz__zz_shift_dataOut_10_1_4,_zz__zz_shift_dataOut_10_1_5};
    end
    if(when_Quan_l130_11) begin
      _zz_shift_dataOut_11_1 <= ($signed(_zz__zz_shift_dataOut_11_1) + $signed(_zz__zz_shift_dataOut_11_1_3));
    end else begin
      _zz_shift_dataOut_11_1 <= {_zz__zz_shift_dataOut_11_1_4,_zz__zz_shift_dataOut_11_1_5};
    end
    if(when_Quan_l130_12) begin
      _zz_shift_dataOut_12_1 <= ($signed(_zz__zz_shift_dataOut_12_1) + $signed(_zz__zz_shift_dataOut_12_1_3));
    end else begin
      _zz_shift_dataOut_12_1 <= {_zz__zz_shift_dataOut_12_1_4,_zz__zz_shift_dataOut_12_1_5};
    end
    if(when_Quan_l130_13) begin
      _zz_shift_dataOut_13_1 <= ($signed(_zz__zz_shift_dataOut_13_1) + $signed(_zz__zz_shift_dataOut_13_1_3));
    end else begin
      _zz_shift_dataOut_13_1 <= {_zz__zz_shift_dataOut_13_1_4,_zz__zz_shift_dataOut_13_1_5};
    end
    if(when_Quan_l130_14) begin
      _zz_shift_dataOut_14_1 <= ($signed(_zz__zz_shift_dataOut_14_1) + $signed(_zz__zz_shift_dataOut_14_1_3));
    end else begin
      _zz_shift_dataOut_14_1 <= {_zz__zz_shift_dataOut_14_1_4,_zz__zz_shift_dataOut_14_1_5};
    end
    if(when_Quan_l130_15) begin
      _zz_shift_dataOut_15_1 <= ($signed(_zz__zz_shift_dataOut_15_1) + $signed(_zz__zz_shift_dataOut_15_1_3));
    end else begin
      _zz_shift_dataOut_15_1 <= {_zz__zz_shift_dataOut_15_1_4,_zz__zz_shift_dataOut_15_1_5};
    end
  end


endmodule

module Scale (
  input      [47:0]   Scale_dataIn_0,
  input      [47:0]   Scale_dataIn_1,
  input      [47:0]   Scale_dataIn_2,
  input      [47:0]   Scale_dataIn_3,
  input      [47:0]   Scale_dataIn_4,
  input      [47:0]   Scale_dataIn_5,
  input      [47:0]   Scale_dataIn_6,
  input      [47:0]   Scale_dataIn_7,
  input      [47:0]   Scale_dataIn_8,
  input      [47:0]   Scale_dataIn_9,
  input      [47:0]   Scale_dataIn_10,
  input      [47:0]   Scale_dataIn_11,
  input      [47:0]   Scale_dataIn_12,
  input      [47:0]   Scale_dataIn_13,
  input      [47:0]   Scale_dataIn_14,
  input      [47:0]   Scale_dataIn_15,
  input      [31:0]   Scale_quan_0,
  input      [31:0]   Scale_quan_1,
  input      [31:0]   Scale_quan_2,
  input      [31:0]   Scale_quan_3,
  input      [31:0]   Scale_quan_4,
  input      [31:0]   Scale_quan_5,
  input      [31:0]   Scale_quan_6,
  input      [31:0]   Scale_quan_7,
  input      [31:0]   Scale_quan_8,
  input      [31:0]   Scale_quan_9,
  input      [31:0]   Scale_quan_10,
  input      [31:0]   Scale_quan_11,
  input      [31:0]   Scale_quan_12,
  input      [31:0]   Scale_quan_13,
  input      [31:0]   Scale_quan_14,
  input      [31:0]   Scale_quan_15,
  output     [31:0]   Scale_dataOut_0,
  output     [31:0]   Scale_dataOut_1,
  output     [31:0]   Scale_dataOut_2,
  output     [31:0]   Scale_dataOut_3,
  output     [31:0]   Scale_dataOut_4,
  output     [31:0]   Scale_dataOut_5,
  output     [31:0]   Scale_dataOut_6,
  output     [31:0]   Scale_dataOut_7,
  output     [31:0]   Scale_dataOut_8,
  output     [31:0]   Scale_dataOut_9,
  output     [31:0]   Scale_dataOut_10,
  output     [31:0]   Scale_dataOut_11,
  output     [31:0]   Scale_dataOut_12,
  output     [31:0]   Scale_dataOut_13,
  output     [31:0]   Scale_dataOut_14,
  output     [31:0]   Scale_dataOut_15,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [31:0]   mul_P;
  wire       [31:0]   mul_1_P;
  wire       [31:0]   mul_2_P;
  wire       [31:0]   mul_3_P;
  wire       [31:0]   mul_4_P;
  wire       [31:0]   mul_5_P;
  wire       [31:0]   mul_6_P;
  wire       [31:0]   mul_7_P;
  wire       [31:0]   mul_8_P;
  wire       [31:0]   mul_9_P;
  wire       [31:0]   mul_10_P;
  wire       [31:0]   mul_11_P;
  wire       [31:0]   mul_12_P;
  wire       [31:0]   mul_13_P;
  wire       [31:0]   mul_14_P;
  wire       [31:0]   mul_15_P;
  wire       [31:0]   scaleMulOut_0;
  wire       [31:0]   scaleMulOut_1;
  wire       [31:0]   scaleMulOut_2;
  wire       [31:0]   scaleMulOut_3;
  wire       [31:0]   scaleMulOut_4;
  wire       [31:0]   scaleMulOut_5;
  wire       [31:0]   scaleMulOut_6;
  wire       [31:0]   scaleMulOut_7;
  wire       [31:0]   scaleMulOut_8;
  wire       [31:0]   scaleMulOut_9;
  wire       [31:0]   scaleMulOut_10;
  wire       [31:0]   scaleMulOut_11;
  wire       [31:0]   scaleMulOut_12;
  wire       [31:0]   scaleMulOut_13;
  wire       [31:0]   scaleMulOut_14;
  wire       [31:0]   scaleMulOut_15;
  reg        [31:0]   scaleMulOut_0_regNext;
  reg        [31:0]   scaleMulOut_1_regNext;
  reg        [31:0]   scaleMulOut_2_regNext;
  reg        [31:0]   scaleMulOut_3_regNext;
  reg        [31:0]   scaleMulOut_4_regNext;
  reg        [31:0]   scaleMulOut_5_regNext;
  reg        [31:0]   scaleMulOut_6_regNext;
  reg        [31:0]   scaleMulOut_7_regNext;
  reg        [31:0]   scaleMulOut_8_regNext;
  reg        [31:0]   scaleMulOut_9_regNext;
  reg        [31:0]   scaleMulOut_10_regNext;
  reg        [31:0]   scaleMulOut_11_regNext;
  reg        [31:0]   scaleMulOut_12_regNext;
  reg        [31:0]   scaleMulOut_13_regNext;
  reg        [31:0]   scaleMulOut_14_regNext;
  reg        [31:0]   scaleMulOut_15_regNext;

  scaleMul mul (
    .A   (Scale_dataIn_0[47:0]), //i
    .B   (Scale_quan_0[31:0]  ), //i
    .P   (mul_P[31:0]         ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_1 (
    .A   (Scale_dataIn_1[47:0]), //i
    .B   (Scale_quan_1[31:0]  ), //i
    .P   (mul_1_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_2 (
    .A   (Scale_dataIn_2[47:0]), //i
    .B   (Scale_quan_2[31:0]  ), //i
    .P   (mul_2_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_3 (
    .A   (Scale_dataIn_3[47:0]), //i
    .B   (Scale_quan_3[31:0]  ), //i
    .P   (mul_3_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_4 (
    .A   (Scale_dataIn_4[47:0]), //i
    .B   (Scale_quan_4[31:0]  ), //i
    .P   (mul_4_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_5 (
    .A   (Scale_dataIn_5[47:0]), //i
    .B   (Scale_quan_5[31:0]  ), //i
    .P   (mul_5_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_6 (
    .A   (Scale_dataIn_6[47:0]), //i
    .B   (Scale_quan_6[31:0]  ), //i
    .P   (mul_6_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_7 (
    .A   (Scale_dataIn_7[47:0]), //i
    .B   (Scale_quan_7[31:0]  ), //i
    .P   (mul_7_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_8 (
    .A   (Scale_dataIn_8[47:0]), //i
    .B   (Scale_quan_8[31:0]  ), //i
    .P   (mul_8_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_9 (
    .A   (Scale_dataIn_9[47:0]), //i
    .B   (Scale_quan_9[31:0]  ), //i
    .P   (mul_9_P[31:0]       ), //o
    .CLK (clk                 )  //i
  );
  scaleMul mul_10 (
    .A   (Scale_dataIn_10[47:0]), //i
    .B   (Scale_quan_10[31:0]  ), //i
    .P   (mul_10_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  scaleMul mul_11 (
    .A   (Scale_dataIn_11[47:0]), //i
    .B   (Scale_quan_11[31:0]  ), //i
    .P   (mul_11_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  scaleMul mul_12 (
    .A   (Scale_dataIn_12[47:0]), //i
    .B   (Scale_quan_12[31:0]  ), //i
    .P   (mul_12_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  scaleMul mul_13 (
    .A   (Scale_dataIn_13[47:0]), //i
    .B   (Scale_quan_13[31:0]  ), //i
    .P   (mul_13_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  scaleMul mul_14 (
    .A   (Scale_dataIn_14[47:0]), //i
    .B   (Scale_quan_14[31:0]  ), //i
    .P   (mul_14_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  scaleMul mul_15 (
    .A   (Scale_dataIn_15[47:0]), //i
    .B   (Scale_quan_15[31:0]  ), //i
    .P   (mul_15_P[31:0]       ), //o
    .CLK (clk                  )  //i
  );
  assign scaleMulOut_0 = mul_P;
  assign scaleMulOut_1 = mul_1_P;
  assign scaleMulOut_2 = mul_2_P;
  assign scaleMulOut_3 = mul_3_P;
  assign scaleMulOut_4 = mul_4_P;
  assign scaleMulOut_5 = mul_5_P;
  assign scaleMulOut_6 = mul_6_P;
  assign scaleMulOut_7 = mul_7_P;
  assign scaleMulOut_8 = mul_8_P;
  assign scaleMulOut_9 = mul_9_P;
  assign scaleMulOut_10 = mul_10_P;
  assign scaleMulOut_11 = mul_11_P;
  assign scaleMulOut_12 = mul_12_P;
  assign scaleMulOut_13 = mul_13_P;
  assign scaleMulOut_14 = mul_14_P;
  assign scaleMulOut_15 = mul_15_P;
  assign Scale_dataOut_0 = scaleMulOut_0_regNext;
  assign Scale_dataOut_1 = scaleMulOut_1_regNext;
  assign Scale_dataOut_2 = scaleMulOut_2_regNext;
  assign Scale_dataOut_3 = scaleMulOut_3_regNext;
  assign Scale_dataOut_4 = scaleMulOut_4_regNext;
  assign Scale_dataOut_5 = scaleMulOut_5_regNext;
  assign Scale_dataOut_6 = scaleMulOut_6_regNext;
  assign Scale_dataOut_7 = scaleMulOut_7_regNext;
  assign Scale_dataOut_8 = scaleMulOut_8_regNext;
  assign Scale_dataOut_9 = scaleMulOut_9_regNext;
  assign Scale_dataOut_10 = scaleMulOut_10_regNext;
  assign Scale_dataOut_11 = scaleMulOut_11_regNext;
  assign Scale_dataOut_12 = scaleMulOut_12_regNext;
  assign Scale_dataOut_13 = scaleMulOut_13_regNext;
  assign Scale_dataOut_14 = scaleMulOut_14_regNext;
  assign Scale_dataOut_15 = scaleMulOut_15_regNext;
  always @(posedge clk) begin
    scaleMulOut_0_regNext <= scaleMulOut_0;
    scaleMulOut_1_regNext <= scaleMulOut_1;
    scaleMulOut_2_regNext <= scaleMulOut_2;
    scaleMulOut_3_regNext <= scaleMulOut_3;
    scaleMulOut_4_regNext <= scaleMulOut_4;
    scaleMulOut_5_regNext <= scaleMulOut_5;
    scaleMulOut_6_regNext <= scaleMulOut_6;
    scaleMulOut_7_regNext <= scaleMulOut_7;
    scaleMulOut_8_regNext <= scaleMulOut_8;
    scaleMulOut_9_regNext <= scaleMulOut_9;
    scaleMulOut_10_regNext <= scaleMulOut_10;
    scaleMulOut_11_regNext <= scaleMulOut_11;
    scaleMulOut_12_regNext <= scaleMulOut_12;
    scaleMulOut_13_regNext <= scaleMulOut_13;
    scaleMulOut_14_regNext <= scaleMulOut_14;
    scaleMulOut_15_regNext <= scaleMulOut_15;
  end


endmodule

module Bias (
  input      [31:0]   Bias_dataIn_0,
  input      [31:0]   Bias_dataIn_1,
  input      [31:0]   Bias_dataIn_2,
  input      [31:0]   Bias_dataIn_3,
  input      [31:0]   Bias_dataIn_4,
  input      [31:0]   Bias_dataIn_5,
  input      [31:0]   Bias_dataIn_6,
  input      [31:0]   Bias_dataIn_7,
  input      [31:0]   Bias_dataIn_8,
  input      [31:0]   Bias_dataIn_9,
  input      [31:0]   Bias_dataIn_10,
  input      [31:0]   Bias_dataIn_11,
  input      [31:0]   Bias_dataIn_12,
  input      [31:0]   Bias_dataIn_13,
  input      [31:0]   Bias_dataIn_14,
  input      [31:0]   Bias_dataIn_15,
  input      [31:0]   Bias_quan_0,
  input      [31:0]   Bias_quan_1,
  input      [31:0]   Bias_quan_2,
  input      [31:0]   Bias_quan_3,
  input      [31:0]   Bias_quan_4,
  input      [31:0]   Bias_quan_5,
  input      [31:0]   Bias_quan_6,
  input      [31:0]   Bias_quan_7,
  input      [31:0]   Bias_quan_8,
  input      [31:0]   Bias_quan_9,
  input      [31:0]   Bias_quan_10,
  input      [31:0]   Bias_quan_11,
  input      [31:0]   Bias_quan_12,
  input      [31:0]   Bias_quan_13,
  input      [31:0]   Bias_quan_14,
  input      [31:0]   Bias_quan_15,
  output     [47:0]   Bias_dataOut_0,
  output     [47:0]   Bias_dataOut_1,
  output     [47:0]   Bias_dataOut_2,
  output     [47:0]   Bias_dataOut_3,
  output     [47:0]   Bias_dataOut_4,
  output     [47:0]   Bias_dataOut_5,
  output     [47:0]   Bias_dataOut_6,
  output     [47:0]   Bias_dataOut_7,
  output     [47:0]   Bias_dataOut_8,
  output     [47:0]   Bias_dataOut_9,
  output     [47:0]   Bias_dataOut_10,
  output     [47:0]   Bias_dataOut_11,
  output     [47:0]   Bias_dataOut_12,
  output     [47:0]   Bias_dataOut_13,
  output     [47:0]   Bias_dataOut_14,
  output     [47:0]   Bias_dataOut_15,
  input               clk,
  input               reset,
  input               softReset
);

  wire       [47:0]   addSub_S;
  wire       [47:0]   addSub_1_S;
  wire       [47:0]   addSub_2_S;
  wire       [47:0]   addSub_3_S;
  wire       [47:0]   addSub_4_S;
  wire       [47:0]   addSub_5_S;
  wire       [47:0]   addSub_6_S;
  wire       [47:0]   addSub_7_S;
  wire       [47:0]   addSub_8_S;
  wire       [47:0]   addSub_9_S;
  wire       [47:0]   addSub_10_S;
  wire       [47:0]   addSub_11_S;
  wire       [47:0]   addSub_12_S;
  wire       [47:0]   addSub_13_S;
  wire       [47:0]   addSub_14_S;
  wire       [47:0]   addSub_15_S;
  wire       [15:0]   _zz_dataInTemp_0;
  wire       [7:0]    _zz_biasInTemp_0;
  wire       [0:0]    _zz_biasInTemp_0_1;
  wire       [8:0]    _zz_biasInTemp_0_2;
  wire       [0:0]    _zz_biasInTemp_0_3;
  wire       [9:0]    _zz_biasInTemp_0_4;
  wire       [0:0]    _zz_biasInTemp_0_5;
  wire       [10:0]   _zz_biasInTemp_0_6;
  wire       [0:0]    _zz_biasInTemp_0_7;
  wire       [11:0]   _zz_biasInTemp_0_8;
  wire       [0:0]    _zz_biasInTemp_0_9;
  wire       [12:0]   _zz_biasInTemp_0_10;
  wire       [0:0]    _zz_biasInTemp_0_11;
  wire       [13:0]   _zz_biasInTemp_0_12;
  wire       [0:0]    _zz_biasInTemp_0_13;
  wire       [14:0]   _zz_biasInTemp_0_14;
  wire       [0:0]    _zz_biasInTemp_0_15;
  wire       [15:0]   _zz_biasInTemp_0_16;
  wire       [0:0]    _zz_biasInTemp_0_17;
  wire       [16:0]   _zz_biasInTemp_0_18;
  wire       [0:0]    _zz_biasInTemp_0_19;
  wire       [17:0]   _zz_biasInTemp_0_20;
  wire       [0:0]    _zz_biasInTemp_0_21;
  wire       [18:0]   _zz_biasInTemp_0_22;
  wire       [0:0]    _zz_biasInTemp_0_23;
  wire       [19:0]   _zz_biasInTemp_0_24;
  wire       [0:0]    _zz_biasInTemp_0_25;
  wire       [20:0]   _zz_biasInTemp_0_26;
  wire       [0:0]    _zz_biasInTemp_0_27;
  wire       [21:0]   _zz_biasInTemp_0_28;
  wire       [0:0]    _zz_biasInTemp_0_29;
  wire       [22:0]   _zz_biasInTemp_0_30;
  wire       [0:0]    _zz_biasInTemp_0_31;
  wire       [23:0]   _zz_biasInTemp_0_32;
  wire       [0:0]    _zz_biasInTemp_0_33;
  wire       [15:0]   _zz_dataInTemp_1;
  wire       [7:0]    _zz_biasInTemp_1;
  wire       [0:0]    _zz_biasInTemp_1_1;
  wire       [8:0]    _zz_biasInTemp_1_2;
  wire       [0:0]    _zz_biasInTemp_1_3;
  wire       [9:0]    _zz_biasInTemp_1_4;
  wire       [0:0]    _zz_biasInTemp_1_5;
  wire       [10:0]   _zz_biasInTemp_1_6;
  wire       [0:0]    _zz_biasInTemp_1_7;
  wire       [11:0]   _zz_biasInTemp_1_8;
  wire       [0:0]    _zz_biasInTemp_1_9;
  wire       [12:0]   _zz_biasInTemp_1_10;
  wire       [0:0]    _zz_biasInTemp_1_11;
  wire       [13:0]   _zz_biasInTemp_1_12;
  wire       [0:0]    _zz_biasInTemp_1_13;
  wire       [14:0]   _zz_biasInTemp_1_14;
  wire       [0:0]    _zz_biasInTemp_1_15;
  wire       [15:0]   _zz_biasInTemp_1_16;
  wire       [0:0]    _zz_biasInTemp_1_17;
  wire       [16:0]   _zz_biasInTemp_1_18;
  wire       [0:0]    _zz_biasInTemp_1_19;
  wire       [17:0]   _zz_biasInTemp_1_20;
  wire       [0:0]    _zz_biasInTemp_1_21;
  wire       [18:0]   _zz_biasInTemp_1_22;
  wire       [0:0]    _zz_biasInTemp_1_23;
  wire       [19:0]   _zz_biasInTemp_1_24;
  wire       [0:0]    _zz_biasInTemp_1_25;
  wire       [20:0]   _zz_biasInTemp_1_26;
  wire       [0:0]    _zz_biasInTemp_1_27;
  wire       [21:0]   _zz_biasInTemp_1_28;
  wire       [0:0]    _zz_biasInTemp_1_29;
  wire       [22:0]   _zz_biasInTemp_1_30;
  wire       [0:0]    _zz_biasInTemp_1_31;
  wire       [23:0]   _zz_biasInTemp_1_32;
  wire       [0:0]    _zz_biasInTemp_1_33;
  wire       [15:0]   _zz_dataInTemp_2;
  wire       [7:0]    _zz_biasInTemp_2;
  wire       [0:0]    _zz_biasInTemp_2_1;
  wire       [8:0]    _zz_biasInTemp_2_2;
  wire       [0:0]    _zz_biasInTemp_2_3;
  wire       [9:0]    _zz_biasInTemp_2_4;
  wire       [0:0]    _zz_biasInTemp_2_5;
  wire       [10:0]   _zz_biasInTemp_2_6;
  wire       [0:0]    _zz_biasInTemp_2_7;
  wire       [11:0]   _zz_biasInTemp_2_8;
  wire       [0:0]    _zz_biasInTemp_2_9;
  wire       [12:0]   _zz_biasInTemp_2_10;
  wire       [0:0]    _zz_biasInTemp_2_11;
  wire       [13:0]   _zz_biasInTemp_2_12;
  wire       [0:0]    _zz_biasInTemp_2_13;
  wire       [14:0]   _zz_biasInTemp_2_14;
  wire       [0:0]    _zz_biasInTemp_2_15;
  wire       [15:0]   _zz_biasInTemp_2_16;
  wire       [0:0]    _zz_biasInTemp_2_17;
  wire       [16:0]   _zz_biasInTemp_2_18;
  wire       [0:0]    _zz_biasInTemp_2_19;
  wire       [17:0]   _zz_biasInTemp_2_20;
  wire       [0:0]    _zz_biasInTemp_2_21;
  wire       [18:0]   _zz_biasInTemp_2_22;
  wire       [0:0]    _zz_biasInTemp_2_23;
  wire       [19:0]   _zz_biasInTemp_2_24;
  wire       [0:0]    _zz_biasInTemp_2_25;
  wire       [20:0]   _zz_biasInTemp_2_26;
  wire       [0:0]    _zz_biasInTemp_2_27;
  wire       [21:0]   _zz_biasInTemp_2_28;
  wire       [0:0]    _zz_biasInTemp_2_29;
  wire       [22:0]   _zz_biasInTemp_2_30;
  wire       [0:0]    _zz_biasInTemp_2_31;
  wire       [23:0]   _zz_biasInTemp_2_32;
  wire       [0:0]    _zz_biasInTemp_2_33;
  wire       [15:0]   _zz_dataInTemp_3;
  wire       [7:0]    _zz_biasInTemp_3;
  wire       [0:0]    _zz_biasInTemp_3_1;
  wire       [8:0]    _zz_biasInTemp_3_2;
  wire       [0:0]    _zz_biasInTemp_3_3;
  wire       [9:0]    _zz_biasInTemp_3_4;
  wire       [0:0]    _zz_biasInTemp_3_5;
  wire       [10:0]   _zz_biasInTemp_3_6;
  wire       [0:0]    _zz_biasInTemp_3_7;
  wire       [11:0]   _zz_biasInTemp_3_8;
  wire       [0:0]    _zz_biasInTemp_3_9;
  wire       [12:0]   _zz_biasInTemp_3_10;
  wire       [0:0]    _zz_biasInTemp_3_11;
  wire       [13:0]   _zz_biasInTemp_3_12;
  wire       [0:0]    _zz_biasInTemp_3_13;
  wire       [14:0]   _zz_biasInTemp_3_14;
  wire       [0:0]    _zz_biasInTemp_3_15;
  wire       [15:0]   _zz_biasInTemp_3_16;
  wire       [0:0]    _zz_biasInTemp_3_17;
  wire       [16:0]   _zz_biasInTemp_3_18;
  wire       [0:0]    _zz_biasInTemp_3_19;
  wire       [17:0]   _zz_biasInTemp_3_20;
  wire       [0:0]    _zz_biasInTemp_3_21;
  wire       [18:0]   _zz_biasInTemp_3_22;
  wire       [0:0]    _zz_biasInTemp_3_23;
  wire       [19:0]   _zz_biasInTemp_3_24;
  wire       [0:0]    _zz_biasInTemp_3_25;
  wire       [20:0]   _zz_biasInTemp_3_26;
  wire       [0:0]    _zz_biasInTemp_3_27;
  wire       [21:0]   _zz_biasInTemp_3_28;
  wire       [0:0]    _zz_biasInTemp_3_29;
  wire       [22:0]   _zz_biasInTemp_3_30;
  wire       [0:0]    _zz_biasInTemp_3_31;
  wire       [23:0]   _zz_biasInTemp_3_32;
  wire       [0:0]    _zz_biasInTemp_3_33;
  wire       [15:0]   _zz_dataInTemp_4;
  wire       [7:0]    _zz_biasInTemp_4;
  wire       [0:0]    _zz_biasInTemp_4_1;
  wire       [8:0]    _zz_biasInTemp_4_2;
  wire       [0:0]    _zz_biasInTemp_4_3;
  wire       [9:0]    _zz_biasInTemp_4_4;
  wire       [0:0]    _zz_biasInTemp_4_5;
  wire       [10:0]   _zz_biasInTemp_4_6;
  wire       [0:0]    _zz_biasInTemp_4_7;
  wire       [11:0]   _zz_biasInTemp_4_8;
  wire       [0:0]    _zz_biasInTemp_4_9;
  wire       [12:0]   _zz_biasInTemp_4_10;
  wire       [0:0]    _zz_biasInTemp_4_11;
  wire       [13:0]   _zz_biasInTemp_4_12;
  wire       [0:0]    _zz_biasInTemp_4_13;
  wire       [14:0]   _zz_biasInTemp_4_14;
  wire       [0:0]    _zz_biasInTemp_4_15;
  wire       [15:0]   _zz_biasInTemp_4_16;
  wire       [0:0]    _zz_biasInTemp_4_17;
  wire       [16:0]   _zz_biasInTemp_4_18;
  wire       [0:0]    _zz_biasInTemp_4_19;
  wire       [17:0]   _zz_biasInTemp_4_20;
  wire       [0:0]    _zz_biasInTemp_4_21;
  wire       [18:0]   _zz_biasInTemp_4_22;
  wire       [0:0]    _zz_biasInTemp_4_23;
  wire       [19:0]   _zz_biasInTemp_4_24;
  wire       [0:0]    _zz_biasInTemp_4_25;
  wire       [20:0]   _zz_biasInTemp_4_26;
  wire       [0:0]    _zz_biasInTemp_4_27;
  wire       [21:0]   _zz_biasInTemp_4_28;
  wire       [0:0]    _zz_biasInTemp_4_29;
  wire       [22:0]   _zz_biasInTemp_4_30;
  wire       [0:0]    _zz_biasInTemp_4_31;
  wire       [23:0]   _zz_biasInTemp_4_32;
  wire       [0:0]    _zz_biasInTemp_4_33;
  wire       [15:0]   _zz_dataInTemp_5;
  wire       [7:0]    _zz_biasInTemp_5;
  wire       [0:0]    _zz_biasInTemp_5_1;
  wire       [8:0]    _zz_biasInTemp_5_2;
  wire       [0:0]    _zz_biasInTemp_5_3;
  wire       [9:0]    _zz_biasInTemp_5_4;
  wire       [0:0]    _zz_biasInTemp_5_5;
  wire       [10:0]   _zz_biasInTemp_5_6;
  wire       [0:0]    _zz_biasInTemp_5_7;
  wire       [11:0]   _zz_biasInTemp_5_8;
  wire       [0:0]    _zz_biasInTemp_5_9;
  wire       [12:0]   _zz_biasInTemp_5_10;
  wire       [0:0]    _zz_biasInTemp_5_11;
  wire       [13:0]   _zz_biasInTemp_5_12;
  wire       [0:0]    _zz_biasInTemp_5_13;
  wire       [14:0]   _zz_biasInTemp_5_14;
  wire       [0:0]    _zz_biasInTemp_5_15;
  wire       [15:0]   _zz_biasInTemp_5_16;
  wire       [0:0]    _zz_biasInTemp_5_17;
  wire       [16:0]   _zz_biasInTemp_5_18;
  wire       [0:0]    _zz_biasInTemp_5_19;
  wire       [17:0]   _zz_biasInTemp_5_20;
  wire       [0:0]    _zz_biasInTemp_5_21;
  wire       [18:0]   _zz_biasInTemp_5_22;
  wire       [0:0]    _zz_biasInTemp_5_23;
  wire       [19:0]   _zz_biasInTemp_5_24;
  wire       [0:0]    _zz_biasInTemp_5_25;
  wire       [20:0]   _zz_biasInTemp_5_26;
  wire       [0:0]    _zz_biasInTemp_5_27;
  wire       [21:0]   _zz_biasInTemp_5_28;
  wire       [0:0]    _zz_biasInTemp_5_29;
  wire       [22:0]   _zz_biasInTemp_5_30;
  wire       [0:0]    _zz_biasInTemp_5_31;
  wire       [23:0]   _zz_biasInTemp_5_32;
  wire       [0:0]    _zz_biasInTemp_5_33;
  wire       [15:0]   _zz_dataInTemp_6;
  wire       [7:0]    _zz_biasInTemp_6;
  wire       [0:0]    _zz_biasInTemp_6_1;
  wire       [8:0]    _zz_biasInTemp_6_2;
  wire       [0:0]    _zz_biasInTemp_6_3;
  wire       [9:0]    _zz_biasInTemp_6_4;
  wire       [0:0]    _zz_biasInTemp_6_5;
  wire       [10:0]   _zz_biasInTemp_6_6;
  wire       [0:0]    _zz_biasInTemp_6_7;
  wire       [11:0]   _zz_biasInTemp_6_8;
  wire       [0:0]    _zz_biasInTemp_6_9;
  wire       [12:0]   _zz_biasInTemp_6_10;
  wire       [0:0]    _zz_biasInTemp_6_11;
  wire       [13:0]   _zz_biasInTemp_6_12;
  wire       [0:0]    _zz_biasInTemp_6_13;
  wire       [14:0]   _zz_biasInTemp_6_14;
  wire       [0:0]    _zz_biasInTemp_6_15;
  wire       [15:0]   _zz_biasInTemp_6_16;
  wire       [0:0]    _zz_biasInTemp_6_17;
  wire       [16:0]   _zz_biasInTemp_6_18;
  wire       [0:0]    _zz_biasInTemp_6_19;
  wire       [17:0]   _zz_biasInTemp_6_20;
  wire       [0:0]    _zz_biasInTemp_6_21;
  wire       [18:0]   _zz_biasInTemp_6_22;
  wire       [0:0]    _zz_biasInTemp_6_23;
  wire       [19:0]   _zz_biasInTemp_6_24;
  wire       [0:0]    _zz_biasInTemp_6_25;
  wire       [20:0]   _zz_biasInTemp_6_26;
  wire       [0:0]    _zz_biasInTemp_6_27;
  wire       [21:0]   _zz_biasInTemp_6_28;
  wire       [0:0]    _zz_biasInTemp_6_29;
  wire       [22:0]   _zz_biasInTemp_6_30;
  wire       [0:0]    _zz_biasInTemp_6_31;
  wire       [23:0]   _zz_biasInTemp_6_32;
  wire       [0:0]    _zz_biasInTemp_6_33;
  wire       [15:0]   _zz_dataInTemp_7;
  wire       [7:0]    _zz_biasInTemp_7;
  wire       [0:0]    _zz_biasInTemp_7_1;
  wire       [8:0]    _zz_biasInTemp_7_2;
  wire       [0:0]    _zz_biasInTemp_7_3;
  wire       [9:0]    _zz_biasInTemp_7_4;
  wire       [0:0]    _zz_biasInTemp_7_5;
  wire       [10:0]   _zz_biasInTemp_7_6;
  wire       [0:0]    _zz_biasInTemp_7_7;
  wire       [11:0]   _zz_biasInTemp_7_8;
  wire       [0:0]    _zz_biasInTemp_7_9;
  wire       [12:0]   _zz_biasInTemp_7_10;
  wire       [0:0]    _zz_biasInTemp_7_11;
  wire       [13:0]   _zz_biasInTemp_7_12;
  wire       [0:0]    _zz_biasInTemp_7_13;
  wire       [14:0]   _zz_biasInTemp_7_14;
  wire       [0:0]    _zz_biasInTemp_7_15;
  wire       [15:0]   _zz_biasInTemp_7_16;
  wire       [0:0]    _zz_biasInTemp_7_17;
  wire       [16:0]   _zz_biasInTemp_7_18;
  wire       [0:0]    _zz_biasInTemp_7_19;
  wire       [17:0]   _zz_biasInTemp_7_20;
  wire       [0:0]    _zz_biasInTemp_7_21;
  wire       [18:0]   _zz_biasInTemp_7_22;
  wire       [0:0]    _zz_biasInTemp_7_23;
  wire       [19:0]   _zz_biasInTemp_7_24;
  wire       [0:0]    _zz_biasInTemp_7_25;
  wire       [20:0]   _zz_biasInTemp_7_26;
  wire       [0:0]    _zz_biasInTemp_7_27;
  wire       [21:0]   _zz_biasInTemp_7_28;
  wire       [0:0]    _zz_biasInTemp_7_29;
  wire       [22:0]   _zz_biasInTemp_7_30;
  wire       [0:0]    _zz_biasInTemp_7_31;
  wire       [23:0]   _zz_biasInTemp_7_32;
  wire       [0:0]    _zz_biasInTemp_7_33;
  wire       [15:0]   _zz_dataInTemp_8;
  wire       [7:0]    _zz_biasInTemp_8;
  wire       [0:0]    _zz_biasInTemp_8_1;
  wire       [8:0]    _zz_biasInTemp_8_2;
  wire       [0:0]    _zz_biasInTemp_8_3;
  wire       [9:0]    _zz_biasInTemp_8_4;
  wire       [0:0]    _zz_biasInTemp_8_5;
  wire       [10:0]   _zz_biasInTemp_8_6;
  wire       [0:0]    _zz_biasInTemp_8_7;
  wire       [11:0]   _zz_biasInTemp_8_8;
  wire       [0:0]    _zz_biasInTemp_8_9;
  wire       [12:0]   _zz_biasInTemp_8_10;
  wire       [0:0]    _zz_biasInTemp_8_11;
  wire       [13:0]   _zz_biasInTemp_8_12;
  wire       [0:0]    _zz_biasInTemp_8_13;
  wire       [14:0]   _zz_biasInTemp_8_14;
  wire       [0:0]    _zz_biasInTemp_8_15;
  wire       [15:0]   _zz_biasInTemp_8_16;
  wire       [0:0]    _zz_biasInTemp_8_17;
  wire       [16:0]   _zz_biasInTemp_8_18;
  wire       [0:0]    _zz_biasInTemp_8_19;
  wire       [17:0]   _zz_biasInTemp_8_20;
  wire       [0:0]    _zz_biasInTemp_8_21;
  wire       [18:0]   _zz_biasInTemp_8_22;
  wire       [0:0]    _zz_biasInTemp_8_23;
  wire       [19:0]   _zz_biasInTemp_8_24;
  wire       [0:0]    _zz_biasInTemp_8_25;
  wire       [20:0]   _zz_biasInTemp_8_26;
  wire       [0:0]    _zz_biasInTemp_8_27;
  wire       [21:0]   _zz_biasInTemp_8_28;
  wire       [0:0]    _zz_biasInTemp_8_29;
  wire       [22:0]   _zz_biasInTemp_8_30;
  wire       [0:0]    _zz_biasInTemp_8_31;
  wire       [23:0]   _zz_biasInTemp_8_32;
  wire       [0:0]    _zz_biasInTemp_8_33;
  wire       [15:0]   _zz_dataInTemp_9;
  wire       [7:0]    _zz_biasInTemp_9;
  wire       [0:0]    _zz_biasInTemp_9_1;
  wire       [8:0]    _zz_biasInTemp_9_2;
  wire       [0:0]    _zz_biasInTemp_9_3;
  wire       [9:0]    _zz_biasInTemp_9_4;
  wire       [0:0]    _zz_biasInTemp_9_5;
  wire       [10:0]   _zz_biasInTemp_9_6;
  wire       [0:0]    _zz_biasInTemp_9_7;
  wire       [11:0]   _zz_biasInTemp_9_8;
  wire       [0:0]    _zz_biasInTemp_9_9;
  wire       [12:0]   _zz_biasInTemp_9_10;
  wire       [0:0]    _zz_biasInTemp_9_11;
  wire       [13:0]   _zz_biasInTemp_9_12;
  wire       [0:0]    _zz_biasInTemp_9_13;
  wire       [14:0]   _zz_biasInTemp_9_14;
  wire       [0:0]    _zz_biasInTemp_9_15;
  wire       [15:0]   _zz_biasInTemp_9_16;
  wire       [0:0]    _zz_biasInTemp_9_17;
  wire       [16:0]   _zz_biasInTemp_9_18;
  wire       [0:0]    _zz_biasInTemp_9_19;
  wire       [17:0]   _zz_biasInTemp_9_20;
  wire       [0:0]    _zz_biasInTemp_9_21;
  wire       [18:0]   _zz_biasInTemp_9_22;
  wire       [0:0]    _zz_biasInTemp_9_23;
  wire       [19:0]   _zz_biasInTemp_9_24;
  wire       [0:0]    _zz_biasInTemp_9_25;
  wire       [20:0]   _zz_biasInTemp_9_26;
  wire       [0:0]    _zz_biasInTemp_9_27;
  wire       [21:0]   _zz_biasInTemp_9_28;
  wire       [0:0]    _zz_biasInTemp_9_29;
  wire       [22:0]   _zz_biasInTemp_9_30;
  wire       [0:0]    _zz_biasInTemp_9_31;
  wire       [23:0]   _zz_biasInTemp_9_32;
  wire       [0:0]    _zz_biasInTemp_9_33;
  wire       [15:0]   _zz_dataInTemp_10;
  wire       [7:0]    _zz_biasInTemp_10;
  wire       [0:0]    _zz_biasInTemp_10_1;
  wire       [8:0]    _zz_biasInTemp_10_2;
  wire       [0:0]    _zz_biasInTemp_10_3;
  wire       [9:0]    _zz_biasInTemp_10_4;
  wire       [0:0]    _zz_biasInTemp_10_5;
  wire       [10:0]   _zz_biasInTemp_10_6;
  wire       [0:0]    _zz_biasInTemp_10_7;
  wire       [11:0]   _zz_biasInTemp_10_8;
  wire       [0:0]    _zz_biasInTemp_10_9;
  wire       [12:0]   _zz_biasInTemp_10_10;
  wire       [0:0]    _zz_biasInTemp_10_11;
  wire       [13:0]   _zz_biasInTemp_10_12;
  wire       [0:0]    _zz_biasInTemp_10_13;
  wire       [14:0]   _zz_biasInTemp_10_14;
  wire       [0:0]    _zz_biasInTemp_10_15;
  wire       [15:0]   _zz_biasInTemp_10_16;
  wire       [0:0]    _zz_biasInTemp_10_17;
  wire       [16:0]   _zz_biasInTemp_10_18;
  wire       [0:0]    _zz_biasInTemp_10_19;
  wire       [17:0]   _zz_biasInTemp_10_20;
  wire       [0:0]    _zz_biasInTemp_10_21;
  wire       [18:0]   _zz_biasInTemp_10_22;
  wire       [0:0]    _zz_biasInTemp_10_23;
  wire       [19:0]   _zz_biasInTemp_10_24;
  wire       [0:0]    _zz_biasInTemp_10_25;
  wire       [20:0]   _zz_biasInTemp_10_26;
  wire       [0:0]    _zz_biasInTemp_10_27;
  wire       [21:0]   _zz_biasInTemp_10_28;
  wire       [0:0]    _zz_biasInTemp_10_29;
  wire       [22:0]   _zz_biasInTemp_10_30;
  wire       [0:0]    _zz_biasInTemp_10_31;
  wire       [23:0]   _zz_biasInTemp_10_32;
  wire       [0:0]    _zz_biasInTemp_10_33;
  wire       [15:0]   _zz_dataInTemp_11;
  wire       [7:0]    _zz_biasInTemp_11;
  wire       [0:0]    _zz_biasInTemp_11_1;
  wire       [8:0]    _zz_biasInTemp_11_2;
  wire       [0:0]    _zz_biasInTemp_11_3;
  wire       [9:0]    _zz_biasInTemp_11_4;
  wire       [0:0]    _zz_biasInTemp_11_5;
  wire       [10:0]   _zz_biasInTemp_11_6;
  wire       [0:0]    _zz_biasInTemp_11_7;
  wire       [11:0]   _zz_biasInTemp_11_8;
  wire       [0:0]    _zz_biasInTemp_11_9;
  wire       [12:0]   _zz_biasInTemp_11_10;
  wire       [0:0]    _zz_biasInTemp_11_11;
  wire       [13:0]   _zz_biasInTemp_11_12;
  wire       [0:0]    _zz_biasInTemp_11_13;
  wire       [14:0]   _zz_biasInTemp_11_14;
  wire       [0:0]    _zz_biasInTemp_11_15;
  wire       [15:0]   _zz_biasInTemp_11_16;
  wire       [0:0]    _zz_biasInTemp_11_17;
  wire       [16:0]   _zz_biasInTemp_11_18;
  wire       [0:0]    _zz_biasInTemp_11_19;
  wire       [17:0]   _zz_biasInTemp_11_20;
  wire       [0:0]    _zz_biasInTemp_11_21;
  wire       [18:0]   _zz_biasInTemp_11_22;
  wire       [0:0]    _zz_biasInTemp_11_23;
  wire       [19:0]   _zz_biasInTemp_11_24;
  wire       [0:0]    _zz_biasInTemp_11_25;
  wire       [20:0]   _zz_biasInTemp_11_26;
  wire       [0:0]    _zz_biasInTemp_11_27;
  wire       [21:0]   _zz_biasInTemp_11_28;
  wire       [0:0]    _zz_biasInTemp_11_29;
  wire       [22:0]   _zz_biasInTemp_11_30;
  wire       [0:0]    _zz_biasInTemp_11_31;
  wire       [23:0]   _zz_biasInTemp_11_32;
  wire       [0:0]    _zz_biasInTemp_11_33;
  wire       [15:0]   _zz_dataInTemp_12;
  wire       [7:0]    _zz_biasInTemp_12;
  wire       [0:0]    _zz_biasInTemp_12_1;
  wire       [8:0]    _zz_biasInTemp_12_2;
  wire       [0:0]    _zz_biasInTemp_12_3;
  wire       [9:0]    _zz_biasInTemp_12_4;
  wire       [0:0]    _zz_biasInTemp_12_5;
  wire       [10:0]   _zz_biasInTemp_12_6;
  wire       [0:0]    _zz_biasInTemp_12_7;
  wire       [11:0]   _zz_biasInTemp_12_8;
  wire       [0:0]    _zz_biasInTemp_12_9;
  wire       [12:0]   _zz_biasInTemp_12_10;
  wire       [0:0]    _zz_biasInTemp_12_11;
  wire       [13:0]   _zz_biasInTemp_12_12;
  wire       [0:0]    _zz_biasInTemp_12_13;
  wire       [14:0]   _zz_biasInTemp_12_14;
  wire       [0:0]    _zz_biasInTemp_12_15;
  wire       [15:0]   _zz_biasInTemp_12_16;
  wire       [0:0]    _zz_biasInTemp_12_17;
  wire       [16:0]   _zz_biasInTemp_12_18;
  wire       [0:0]    _zz_biasInTemp_12_19;
  wire       [17:0]   _zz_biasInTemp_12_20;
  wire       [0:0]    _zz_biasInTemp_12_21;
  wire       [18:0]   _zz_biasInTemp_12_22;
  wire       [0:0]    _zz_biasInTemp_12_23;
  wire       [19:0]   _zz_biasInTemp_12_24;
  wire       [0:0]    _zz_biasInTemp_12_25;
  wire       [20:0]   _zz_biasInTemp_12_26;
  wire       [0:0]    _zz_biasInTemp_12_27;
  wire       [21:0]   _zz_biasInTemp_12_28;
  wire       [0:0]    _zz_biasInTemp_12_29;
  wire       [22:0]   _zz_biasInTemp_12_30;
  wire       [0:0]    _zz_biasInTemp_12_31;
  wire       [23:0]   _zz_biasInTemp_12_32;
  wire       [0:0]    _zz_biasInTemp_12_33;
  wire       [15:0]   _zz_dataInTemp_13;
  wire       [7:0]    _zz_biasInTemp_13;
  wire       [0:0]    _zz_biasInTemp_13_1;
  wire       [8:0]    _zz_biasInTemp_13_2;
  wire       [0:0]    _zz_biasInTemp_13_3;
  wire       [9:0]    _zz_biasInTemp_13_4;
  wire       [0:0]    _zz_biasInTemp_13_5;
  wire       [10:0]   _zz_biasInTemp_13_6;
  wire       [0:0]    _zz_biasInTemp_13_7;
  wire       [11:0]   _zz_biasInTemp_13_8;
  wire       [0:0]    _zz_biasInTemp_13_9;
  wire       [12:0]   _zz_biasInTemp_13_10;
  wire       [0:0]    _zz_biasInTemp_13_11;
  wire       [13:0]   _zz_biasInTemp_13_12;
  wire       [0:0]    _zz_biasInTemp_13_13;
  wire       [14:0]   _zz_biasInTemp_13_14;
  wire       [0:0]    _zz_biasInTemp_13_15;
  wire       [15:0]   _zz_biasInTemp_13_16;
  wire       [0:0]    _zz_biasInTemp_13_17;
  wire       [16:0]   _zz_biasInTemp_13_18;
  wire       [0:0]    _zz_biasInTemp_13_19;
  wire       [17:0]   _zz_biasInTemp_13_20;
  wire       [0:0]    _zz_biasInTemp_13_21;
  wire       [18:0]   _zz_biasInTemp_13_22;
  wire       [0:0]    _zz_biasInTemp_13_23;
  wire       [19:0]   _zz_biasInTemp_13_24;
  wire       [0:0]    _zz_biasInTemp_13_25;
  wire       [20:0]   _zz_biasInTemp_13_26;
  wire       [0:0]    _zz_biasInTemp_13_27;
  wire       [21:0]   _zz_biasInTemp_13_28;
  wire       [0:0]    _zz_biasInTemp_13_29;
  wire       [22:0]   _zz_biasInTemp_13_30;
  wire       [0:0]    _zz_biasInTemp_13_31;
  wire       [23:0]   _zz_biasInTemp_13_32;
  wire       [0:0]    _zz_biasInTemp_13_33;
  wire       [15:0]   _zz_dataInTemp_14;
  wire       [7:0]    _zz_biasInTemp_14;
  wire       [0:0]    _zz_biasInTemp_14_1;
  wire       [8:0]    _zz_biasInTemp_14_2;
  wire       [0:0]    _zz_biasInTemp_14_3;
  wire       [9:0]    _zz_biasInTemp_14_4;
  wire       [0:0]    _zz_biasInTemp_14_5;
  wire       [10:0]   _zz_biasInTemp_14_6;
  wire       [0:0]    _zz_biasInTemp_14_7;
  wire       [11:0]   _zz_biasInTemp_14_8;
  wire       [0:0]    _zz_biasInTemp_14_9;
  wire       [12:0]   _zz_biasInTemp_14_10;
  wire       [0:0]    _zz_biasInTemp_14_11;
  wire       [13:0]   _zz_biasInTemp_14_12;
  wire       [0:0]    _zz_biasInTemp_14_13;
  wire       [14:0]   _zz_biasInTemp_14_14;
  wire       [0:0]    _zz_biasInTemp_14_15;
  wire       [15:0]   _zz_biasInTemp_14_16;
  wire       [0:0]    _zz_biasInTemp_14_17;
  wire       [16:0]   _zz_biasInTemp_14_18;
  wire       [0:0]    _zz_biasInTemp_14_19;
  wire       [17:0]   _zz_biasInTemp_14_20;
  wire       [0:0]    _zz_biasInTemp_14_21;
  wire       [18:0]   _zz_biasInTemp_14_22;
  wire       [0:0]    _zz_biasInTemp_14_23;
  wire       [19:0]   _zz_biasInTemp_14_24;
  wire       [0:0]    _zz_biasInTemp_14_25;
  wire       [20:0]   _zz_biasInTemp_14_26;
  wire       [0:0]    _zz_biasInTemp_14_27;
  wire       [21:0]   _zz_biasInTemp_14_28;
  wire       [0:0]    _zz_biasInTemp_14_29;
  wire       [22:0]   _zz_biasInTemp_14_30;
  wire       [0:0]    _zz_biasInTemp_14_31;
  wire       [23:0]   _zz_biasInTemp_14_32;
  wire       [0:0]    _zz_biasInTemp_14_33;
  wire       [15:0]   _zz_dataInTemp_15;
  wire       [7:0]    _zz_biasInTemp_15;
  wire       [0:0]    _zz_biasInTemp_15_1;
  wire       [8:0]    _zz_biasInTemp_15_2;
  wire       [0:0]    _zz_biasInTemp_15_3;
  wire       [9:0]    _zz_biasInTemp_15_4;
  wire       [0:0]    _zz_biasInTemp_15_5;
  wire       [10:0]   _zz_biasInTemp_15_6;
  wire       [0:0]    _zz_biasInTemp_15_7;
  wire       [11:0]   _zz_biasInTemp_15_8;
  wire       [0:0]    _zz_biasInTemp_15_9;
  wire       [12:0]   _zz_biasInTemp_15_10;
  wire       [0:0]    _zz_biasInTemp_15_11;
  wire       [13:0]   _zz_biasInTemp_15_12;
  wire       [0:0]    _zz_biasInTemp_15_13;
  wire       [14:0]   _zz_biasInTemp_15_14;
  wire       [0:0]    _zz_biasInTemp_15_15;
  wire       [15:0]   _zz_biasInTemp_15_16;
  wire       [0:0]    _zz_biasInTemp_15_17;
  wire       [16:0]   _zz_biasInTemp_15_18;
  wire       [0:0]    _zz_biasInTemp_15_19;
  wire       [17:0]   _zz_biasInTemp_15_20;
  wire       [0:0]    _zz_biasInTemp_15_21;
  wire       [18:0]   _zz_biasInTemp_15_22;
  wire       [0:0]    _zz_biasInTemp_15_23;
  wire       [19:0]   _zz_biasInTemp_15_24;
  wire       [0:0]    _zz_biasInTemp_15_25;
  wire       [20:0]   _zz_biasInTemp_15_26;
  wire       [0:0]    _zz_biasInTemp_15_27;
  wire       [21:0]   _zz_biasInTemp_15_28;
  wire       [0:0]    _zz_biasInTemp_15_29;
  wire       [22:0]   _zz_biasInTemp_15_30;
  wire       [0:0]    _zz_biasInTemp_15_31;
  wire       [23:0]   _zz_biasInTemp_15_32;
  wire       [0:0]    _zz_biasInTemp_15_33;
  reg        [47:0]   dataInTemp_0;
  reg        [47:0]   dataInTemp_1;
  reg        [47:0]   dataInTemp_2;
  reg        [47:0]   dataInTemp_3;
  reg        [47:0]   dataInTemp_4;
  reg        [47:0]   dataInTemp_5;
  reg        [47:0]   dataInTemp_6;
  reg        [47:0]   dataInTemp_7;
  reg        [47:0]   dataInTemp_8;
  reg        [47:0]   dataInTemp_9;
  reg        [47:0]   dataInTemp_10;
  reg        [47:0]   dataInTemp_11;
  reg        [47:0]   dataInTemp_12;
  reg        [47:0]   dataInTemp_13;
  reg        [47:0]   dataInTemp_14;
  reg        [47:0]   dataInTemp_15;
  reg        [47:0]   biasInTemp_0;
  reg        [47:0]   biasInTemp_1;
  reg        [47:0]   biasInTemp_2;
  reg        [47:0]   biasInTemp_3;
  reg        [47:0]   biasInTemp_4;
  reg        [47:0]   biasInTemp_5;
  reg        [47:0]   biasInTemp_6;
  reg        [47:0]   biasInTemp_7;
  reg        [47:0]   biasInTemp_8;
  reg        [47:0]   biasInTemp_9;
  reg        [47:0]   biasInTemp_10;
  reg        [47:0]   biasInTemp_11;
  reg        [47:0]   biasInTemp_12;
  reg        [47:0]   biasInTemp_13;
  reg        [47:0]   biasInTemp_14;
  reg        [47:0]   biasInTemp_15;
  wire       [6:0]    switch_Quan_l67;
  wire       [6:0]    switch_Quan_l67_1;
  wire       [6:0]    switch_Quan_l67_2;
  wire       [6:0]    switch_Quan_l67_3;
  wire       [6:0]    switch_Quan_l67_4;
  wire       [6:0]    switch_Quan_l67_5;
  wire       [6:0]    switch_Quan_l67_6;
  wire       [6:0]    switch_Quan_l67_7;
  wire       [6:0]    switch_Quan_l67_8;
  wire       [6:0]    switch_Quan_l67_9;
  wire       [6:0]    switch_Quan_l67_10;
  wire       [6:0]    switch_Quan_l67_11;
  wire       [6:0]    switch_Quan_l67_12;
  wire       [6:0]    switch_Quan_l67_13;
  wire       [6:0]    switch_Quan_l67_14;
  wire       [6:0]    switch_Quan_l67_15;

  assign _zz_dataInTemp_0 = 16'h0;
  assign _zz_biasInTemp_0_1 = Bias_quan_0[31];
  assign _zz_biasInTemp_0 = {{7{_zz_biasInTemp_0_1[0]}}, _zz_biasInTemp_0_1};
  assign _zz_biasInTemp_0_3 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_2 = {{8{_zz_biasInTemp_0_3[0]}}, _zz_biasInTemp_0_3};
  assign _zz_biasInTemp_0_5 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_4 = {{9{_zz_biasInTemp_0_5[0]}}, _zz_biasInTemp_0_5};
  assign _zz_biasInTemp_0_7 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_6 = {{10{_zz_biasInTemp_0_7[0]}}, _zz_biasInTemp_0_7};
  assign _zz_biasInTemp_0_9 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_8 = {{11{_zz_biasInTemp_0_9[0]}}, _zz_biasInTemp_0_9};
  assign _zz_biasInTemp_0_11 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_10 = {{12{_zz_biasInTemp_0_11[0]}}, _zz_biasInTemp_0_11};
  assign _zz_biasInTemp_0_13 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_12 = {{13{_zz_biasInTemp_0_13[0]}}, _zz_biasInTemp_0_13};
  assign _zz_biasInTemp_0_15 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_14 = {{14{_zz_biasInTemp_0_15[0]}}, _zz_biasInTemp_0_15};
  assign _zz_biasInTemp_0_17 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_16 = {{15{_zz_biasInTemp_0_17[0]}}, _zz_biasInTemp_0_17};
  assign _zz_biasInTemp_0_19 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_18 = {{16{_zz_biasInTemp_0_19[0]}}, _zz_biasInTemp_0_19};
  assign _zz_biasInTemp_0_21 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_20 = {{17{_zz_biasInTemp_0_21[0]}}, _zz_biasInTemp_0_21};
  assign _zz_biasInTemp_0_23 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_22 = {{18{_zz_biasInTemp_0_23[0]}}, _zz_biasInTemp_0_23};
  assign _zz_biasInTemp_0_25 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_24 = {{19{_zz_biasInTemp_0_25[0]}}, _zz_biasInTemp_0_25};
  assign _zz_biasInTemp_0_27 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_26 = {{20{_zz_biasInTemp_0_27[0]}}, _zz_biasInTemp_0_27};
  assign _zz_biasInTemp_0_29 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_28 = {{21{_zz_biasInTemp_0_29[0]}}, _zz_biasInTemp_0_29};
  assign _zz_biasInTemp_0_31 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_30 = {{22{_zz_biasInTemp_0_31[0]}}, _zz_biasInTemp_0_31};
  assign _zz_biasInTemp_0_33 = Bias_quan_0[31];
  assign _zz_biasInTemp_0_32 = {{23{_zz_biasInTemp_0_33[0]}}, _zz_biasInTemp_0_33};
  assign _zz_dataInTemp_1 = 16'h0;
  assign _zz_biasInTemp_1_1 = Bias_quan_1[31];
  assign _zz_biasInTemp_1 = {{7{_zz_biasInTemp_1_1[0]}}, _zz_biasInTemp_1_1};
  assign _zz_biasInTemp_1_3 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_2 = {{8{_zz_biasInTemp_1_3[0]}}, _zz_biasInTemp_1_3};
  assign _zz_biasInTemp_1_5 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_4 = {{9{_zz_biasInTemp_1_5[0]}}, _zz_biasInTemp_1_5};
  assign _zz_biasInTemp_1_7 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_6 = {{10{_zz_biasInTemp_1_7[0]}}, _zz_biasInTemp_1_7};
  assign _zz_biasInTemp_1_9 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_8 = {{11{_zz_biasInTemp_1_9[0]}}, _zz_biasInTemp_1_9};
  assign _zz_biasInTemp_1_11 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_10 = {{12{_zz_biasInTemp_1_11[0]}}, _zz_biasInTemp_1_11};
  assign _zz_biasInTemp_1_13 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_12 = {{13{_zz_biasInTemp_1_13[0]}}, _zz_biasInTemp_1_13};
  assign _zz_biasInTemp_1_15 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_14 = {{14{_zz_biasInTemp_1_15[0]}}, _zz_biasInTemp_1_15};
  assign _zz_biasInTemp_1_17 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_16 = {{15{_zz_biasInTemp_1_17[0]}}, _zz_biasInTemp_1_17};
  assign _zz_biasInTemp_1_19 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_18 = {{16{_zz_biasInTemp_1_19[0]}}, _zz_biasInTemp_1_19};
  assign _zz_biasInTemp_1_21 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_20 = {{17{_zz_biasInTemp_1_21[0]}}, _zz_biasInTemp_1_21};
  assign _zz_biasInTemp_1_23 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_22 = {{18{_zz_biasInTemp_1_23[0]}}, _zz_biasInTemp_1_23};
  assign _zz_biasInTemp_1_25 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_24 = {{19{_zz_biasInTemp_1_25[0]}}, _zz_biasInTemp_1_25};
  assign _zz_biasInTemp_1_27 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_26 = {{20{_zz_biasInTemp_1_27[0]}}, _zz_biasInTemp_1_27};
  assign _zz_biasInTemp_1_29 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_28 = {{21{_zz_biasInTemp_1_29[0]}}, _zz_biasInTemp_1_29};
  assign _zz_biasInTemp_1_31 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_30 = {{22{_zz_biasInTemp_1_31[0]}}, _zz_biasInTemp_1_31};
  assign _zz_biasInTemp_1_33 = Bias_quan_1[31];
  assign _zz_biasInTemp_1_32 = {{23{_zz_biasInTemp_1_33[0]}}, _zz_biasInTemp_1_33};
  assign _zz_dataInTemp_2 = 16'h0;
  assign _zz_biasInTemp_2_1 = Bias_quan_2[31];
  assign _zz_biasInTemp_2 = {{7{_zz_biasInTemp_2_1[0]}}, _zz_biasInTemp_2_1};
  assign _zz_biasInTemp_2_3 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_2 = {{8{_zz_biasInTemp_2_3[0]}}, _zz_biasInTemp_2_3};
  assign _zz_biasInTemp_2_5 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_4 = {{9{_zz_biasInTemp_2_5[0]}}, _zz_biasInTemp_2_5};
  assign _zz_biasInTemp_2_7 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_6 = {{10{_zz_biasInTemp_2_7[0]}}, _zz_biasInTemp_2_7};
  assign _zz_biasInTemp_2_9 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_8 = {{11{_zz_biasInTemp_2_9[0]}}, _zz_biasInTemp_2_9};
  assign _zz_biasInTemp_2_11 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_10 = {{12{_zz_biasInTemp_2_11[0]}}, _zz_biasInTemp_2_11};
  assign _zz_biasInTemp_2_13 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_12 = {{13{_zz_biasInTemp_2_13[0]}}, _zz_biasInTemp_2_13};
  assign _zz_biasInTemp_2_15 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_14 = {{14{_zz_biasInTemp_2_15[0]}}, _zz_biasInTemp_2_15};
  assign _zz_biasInTemp_2_17 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_16 = {{15{_zz_biasInTemp_2_17[0]}}, _zz_biasInTemp_2_17};
  assign _zz_biasInTemp_2_19 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_18 = {{16{_zz_biasInTemp_2_19[0]}}, _zz_biasInTemp_2_19};
  assign _zz_biasInTemp_2_21 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_20 = {{17{_zz_biasInTemp_2_21[0]}}, _zz_biasInTemp_2_21};
  assign _zz_biasInTemp_2_23 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_22 = {{18{_zz_biasInTemp_2_23[0]}}, _zz_biasInTemp_2_23};
  assign _zz_biasInTemp_2_25 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_24 = {{19{_zz_biasInTemp_2_25[0]}}, _zz_biasInTemp_2_25};
  assign _zz_biasInTemp_2_27 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_26 = {{20{_zz_biasInTemp_2_27[0]}}, _zz_biasInTemp_2_27};
  assign _zz_biasInTemp_2_29 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_28 = {{21{_zz_biasInTemp_2_29[0]}}, _zz_biasInTemp_2_29};
  assign _zz_biasInTemp_2_31 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_30 = {{22{_zz_biasInTemp_2_31[0]}}, _zz_biasInTemp_2_31};
  assign _zz_biasInTemp_2_33 = Bias_quan_2[31];
  assign _zz_biasInTemp_2_32 = {{23{_zz_biasInTemp_2_33[0]}}, _zz_biasInTemp_2_33};
  assign _zz_dataInTemp_3 = 16'h0;
  assign _zz_biasInTemp_3_1 = Bias_quan_3[31];
  assign _zz_biasInTemp_3 = {{7{_zz_biasInTemp_3_1[0]}}, _zz_biasInTemp_3_1};
  assign _zz_biasInTemp_3_3 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_2 = {{8{_zz_biasInTemp_3_3[0]}}, _zz_biasInTemp_3_3};
  assign _zz_biasInTemp_3_5 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_4 = {{9{_zz_biasInTemp_3_5[0]}}, _zz_biasInTemp_3_5};
  assign _zz_biasInTemp_3_7 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_6 = {{10{_zz_biasInTemp_3_7[0]}}, _zz_biasInTemp_3_7};
  assign _zz_biasInTemp_3_9 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_8 = {{11{_zz_biasInTemp_3_9[0]}}, _zz_biasInTemp_3_9};
  assign _zz_biasInTemp_3_11 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_10 = {{12{_zz_biasInTemp_3_11[0]}}, _zz_biasInTemp_3_11};
  assign _zz_biasInTemp_3_13 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_12 = {{13{_zz_biasInTemp_3_13[0]}}, _zz_biasInTemp_3_13};
  assign _zz_biasInTemp_3_15 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_14 = {{14{_zz_biasInTemp_3_15[0]}}, _zz_biasInTemp_3_15};
  assign _zz_biasInTemp_3_17 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_16 = {{15{_zz_biasInTemp_3_17[0]}}, _zz_biasInTemp_3_17};
  assign _zz_biasInTemp_3_19 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_18 = {{16{_zz_biasInTemp_3_19[0]}}, _zz_biasInTemp_3_19};
  assign _zz_biasInTemp_3_21 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_20 = {{17{_zz_biasInTemp_3_21[0]}}, _zz_biasInTemp_3_21};
  assign _zz_biasInTemp_3_23 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_22 = {{18{_zz_biasInTemp_3_23[0]}}, _zz_biasInTemp_3_23};
  assign _zz_biasInTemp_3_25 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_24 = {{19{_zz_biasInTemp_3_25[0]}}, _zz_biasInTemp_3_25};
  assign _zz_biasInTemp_3_27 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_26 = {{20{_zz_biasInTemp_3_27[0]}}, _zz_biasInTemp_3_27};
  assign _zz_biasInTemp_3_29 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_28 = {{21{_zz_biasInTemp_3_29[0]}}, _zz_biasInTemp_3_29};
  assign _zz_biasInTemp_3_31 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_30 = {{22{_zz_biasInTemp_3_31[0]}}, _zz_biasInTemp_3_31};
  assign _zz_biasInTemp_3_33 = Bias_quan_3[31];
  assign _zz_biasInTemp_3_32 = {{23{_zz_biasInTemp_3_33[0]}}, _zz_biasInTemp_3_33};
  assign _zz_dataInTemp_4 = 16'h0;
  assign _zz_biasInTemp_4_1 = Bias_quan_4[31];
  assign _zz_biasInTemp_4 = {{7{_zz_biasInTemp_4_1[0]}}, _zz_biasInTemp_4_1};
  assign _zz_biasInTemp_4_3 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_2 = {{8{_zz_biasInTemp_4_3[0]}}, _zz_biasInTemp_4_3};
  assign _zz_biasInTemp_4_5 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_4 = {{9{_zz_biasInTemp_4_5[0]}}, _zz_biasInTemp_4_5};
  assign _zz_biasInTemp_4_7 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_6 = {{10{_zz_biasInTemp_4_7[0]}}, _zz_biasInTemp_4_7};
  assign _zz_biasInTemp_4_9 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_8 = {{11{_zz_biasInTemp_4_9[0]}}, _zz_biasInTemp_4_9};
  assign _zz_biasInTemp_4_11 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_10 = {{12{_zz_biasInTemp_4_11[0]}}, _zz_biasInTemp_4_11};
  assign _zz_biasInTemp_4_13 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_12 = {{13{_zz_biasInTemp_4_13[0]}}, _zz_biasInTemp_4_13};
  assign _zz_biasInTemp_4_15 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_14 = {{14{_zz_biasInTemp_4_15[0]}}, _zz_biasInTemp_4_15};
  assign _zz_biasInTemp_4_17 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_16 = {{15{_zz_biasInTemp_4_17[0]}}, _zz_biasInTemp_4_17};
  assign _zz_biasInTemp_4_19 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_18 = {{16{_zz_biasInTemp_4_19[0]}}, _zz_biasInTemp_4_19};
  assign _zz_biasInTemp_4_21 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_20 = {{17{_zz_biasInTemp_4_21[0]}}, _zz_biasInTemp_4_21};
  assign _zz_biasInTemp_4_23 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_22 = {{18{_zz_biasInTemp_4_23[0]}}, _zz_biasInTemp_4_23};
  assign _zz_biasInTemp_4_25 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_24 = {{19{_zz_biasInTemp_4_25[0]}}, _zz_biasInTemp_4_25};
  assign _zz_biasInTemp_4_27 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_26 = {{20{_zz_biasInTemp_4_27[0]}}, _zz_biasInTemp_4_27};
  assign _zz_biasInTemp_4_29 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_28 = {{21{_zz_biasInTemp_4_29[0]}}, _zz_biasInTemp_4_29};
  assign _zz_biasInTemp_4_31 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_30 = {{22{_zz_biasInTemp_4_31[0]}}, _zz_biasInTemp_4_31};
  assign _zz_biasInTemp_4_33 = Bias_quan_4[31];
  assign _zz_biasInTemp_4_32 = {{23{_zz_biasInTemp_4_33[0]}}, _zz_biasInTemp_4_33};
  assign _zz_dataInTemp_5 = 16'h0;
  assign _zz_biasInTemp_5_1 = Bias_quan_5[31];
  assign _zz_biasInTemp_5 = {{7{_zz_biasInTemp_5_1[0]}}, _zz_biasInTemp_5_1};
  assign _zz_biasInTemp_5_3 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_2 = {{8{_zz_biasInTemp_5_3[0]}}, _zz_biasInTemp_5_3};
  assign _zz_biasInTemp_5_5 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_4 = {{9{_zz_biasInTemp_5_5[0]}}, _zz_biasInTemp_5_5};
  assign _zz_biasInTemp_5_7 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_6 = {{10{_zz_biasInTemp_5_7[0]}}, _zz_biasInTemp_5_7};
  assign _zz_biasInTemp_5_9 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_8 = {{11{_zz_biasInTemp_5_9[0]}}, _zz_biasInTemp_5_9};
  assign _zz_biasInTemp_5_11 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_10 = {{12{_zz_biasInTemp_5_11[0]}}, _zz_biasInTemp_5_11};
  assign _zz_biasInTemp_5_13 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_12 = {{13{_zz_biasInTemp_5_13[0]}}, _zz_biasInTemp_5_13};
  assign _zz_biasInTemp_5_15 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_14 = {{14{_zz_biasInTemp_5_15[0]}}, _zz_biasInTemp_5_15};
  assign _zz_biasInTemp_5_17 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_16 = {{15{_zz_biasInTemp_5_17[0]}}, _zz_biasInTemp_5_17};
  assign _zz_biasInTemp_5_19 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_18 = {{16{_zz_biasInTemp_5_19[0]}}, _zz_biasInTemp_5_19};
  assign _zz_biasInTemp_5_21 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_20 = {{17{_zz_biasInTemp_5_21[0]}}, _zz_biasInTemp_5_21};
  assign _zz_biasInTemp_5_23 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_22 = {{18{_zz_biasInTemp_5_23[0]}}, _zz_biasInTemp_5_23};
  assign _zz_biasInTemp_5_25 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_24 = {{19{_zz_biasInTemp_5_25[0]}}, _zz_biasInTemp_5_25};
  assign _zz_biasInTemp_5_27 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_26 = {{20{_zz_biasInTemp_5_27[0]}}, _zz_biasInTemp_5_27};
  assign _zz_biasInTemp_5_29 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_28 = {{21{_zz_biasInTemp_5_29[0]}}, _zz_biasInTemp_5_29};
  assign _zz_biasInTemp_5_31 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_30 = {{22{_zz_biasInTemp_5_31[0]}}, _zz_biasInTemp_5_31};
  assign _zz_biasInTemp_5_33 = Bias_quan_5[31];
  assign _zz_biasInTemp_5_32 = {{23{_zz_biasInTemp_5_33[0]}}, _zz_biasInTemp_5_33};
  assign _zz_dataInTemp_6 = 16'h0;
  assign _zz_biasInTemp_6_1 = Bias_quan_6[31];
  assign _zz_biasInTemp_6 = {{7{_zz_biasInTemp_6_1[0]}}, _zz_biasInTemp_6_1};
  assign _zz_biasInTemp_6_3 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_2 = {{8{_zz_biasInTemp_6_3[0]}}, _zz_biasInTemp_6_3};
  assign _zz_biasInTemp_6_5 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_4 = {{9{_zz_biasInTemp_6_5[0]}}, _zz_biasInTemp_6_5};
  assign _zz_biasInTemp_6_7 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_6 = {{10{_zz_biasInTemp_6_7[0]}}, _zz_biasInTemp_6_7};
  assign _zz_biasInTemp_6_9 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_8 = {{11{_zz_biasInTemp_6_9[0]}}, _zz_biasInTemp_6_9};
  assign _zz_biasInTemp_6_11 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_10 = {{12{_zz_biasInTemp_6_11[0]}}, _zz_biasInTemp_6_11};
  assign _zz_biasInTemp_6_13 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_12 = {{13{_zz_biasInTemp_6_13[0]}}, _zz_biasInTemp_6_13};
  assign _zz_biasInTemp_6_15 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_14 = {{14{_zz_biasInTemp_6_15[0]}}, _zz_biasInTemp_6_15};
  assign _zz_biasInTemp_6_17 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_16 = {{15{_zz_biasInTemp_6_17[0]}}, _zz_biasInTemp_6_17};
  assign _zz_biasInTemp_6_19 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_18 = {{16{_zz_biasInTemp_6_19[0]}}, _zz_biasInTemp_6_19};
  assign _zz_biasInTemp_6_21 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_20 = {{17{_zz_biasInTemp_6_21[0]}}, _zz_biasInTemp_6_21};
  assign _zz_biasInTemp_6_23 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_22 = {{18{_zz_biasInTemp_6_23[0]}}, _zz_biasInTemp_6_23};
  assign _zz_biasInTemp_6_25 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_24 = {{19{_zz_biasInTemp_6_25[0]}}, _zz_biasInTemp_6_25};
  assign _zz_biasInTemp_6_27 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_26 = {{20{_zz_biasInTemp_6_27[0]}}, _zz_biasInTemp_6_27};
  assign _zz_biasInTemp_6_29 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_28 = {{21{_zz_biasInTemp_6_29[0]}}, _zz_biasInTemp_6_29};
  assign _zz_biasInTemp_6_31 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_30 = {{22{_zz_biasInTemp_6_31[0]}}, _zz_biasInTemp_6_31};
  assign _zz_biasInTemp_6_33 = Bias_quan_6[31];
  assign _zz_biasInTemp_6_32 = {{23{_zz_biasInTemp_6_33[0]}}, _zz_biasInTemp_6_33};
  assign _zz_dataInTemp_7 = 16'h0;
  assign _zz_biasInTemp_7_1 = Bias_quan_7[31];
  assign _zz_biasInTemp_7 = {{7{_zz_biasInTemp_7_1[0]}}, _zz_biasInTemp_7_1};
  assign _zz_biasInTemp_7_3 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_2 = {{8{_zz_biasInTemp_7_3[0]}}, _zz_biasInTemp_7_3};
  assign _zz_biasInTemp_7_5 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_4 = {{9{_zz_biasInTemp_7_5[0]}}, _zz_biasInTemp_7_5};
  assign _zz_biasInTemp_7_7 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_6 = {{10{_zz_biasInTemp_7_7[0]}}, _zz_biasInTemp_7_7};
  assign _zz_biasInTemp_7_9 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_8 = {{11{_zz_biasInTemp_7_9[0]}}, _zz_biasInTemp_7_9};
  assign _zz_biasInTemp_7_11 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_10 = {{12{_zz_biasInTemp_7_11[0]}}, _zz_biasInTemp_7_11};
  assign _zz_biasInTemp_7_13 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_12 = {{13{_zz_biasInTemp_7_13[0]}}, _zz_biasInTemp_7_13};
  assign _zz_biasInTemp_7_15 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_14 = {{14{_zz_biasInTemp_7_15[0]}}, _zz_biasInTemp_7_15};
  assign _zz_biasInTemp_7_17 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_16 = {{15{_zz_biasInTemp_7_17[0]}}, _zz_biasInTemp_7_17};
  assign _zz_biasInTemp_7_19 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_18 = {{16{_zz_biasInTemp_7_19[0]}}, _zz_biasInTemp_7_19};
  assign _zz_biasInTemp_7_21 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_20 = {{17{_zz_biasInTemp_7_21[0]}}, _zz_biasInTemp_7_21};
  assign _zz_biasInTemp_7_23 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_22 = {{18{_zz_biasInTemp_7_23[0]}}, _zz_biasInTemp_7_23};
  assign _zz_biasInTemp_7_25 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_24 = {{19{_zz_biasInTemp_7_25[0]}}, _zz_biasInTemp_7_25};
  assign _zz_biasInTemp_7_27 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_26 = {{20{_zz_biasInTemp_7_27[0]}}, _zz_biasInTemp_7_27};
  assign _zz_biasInTemp_7_29 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_28 = {{21{_zz_biasInTemp_7_29[0]}}, _zz_biasInTemp_7_29};
  assign _zz_biasInTemp_7_31 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_30 = {{22{_zz_biasInTemp_7_31[0]}}, _zz_biasInTemp_7_31};
  assign _zz_biasInTemp_7_33 = Bias_quan_7[31];
  assign _zz_biasInTemp_7_32 = {{23{_zz_biasInTemp_7_33[0]}}, _zz_biasInTemp_7_33};
  assign _zz_dataInTemp_8 = 16'h0;
  assign _zz_biasInTemp_8_1 = Bias_quan_8[31];
  assign _zz_biasInTemp_8 = {{7{_zz_biasInTemp_8_1[0]}}, _zz_biasInTemp_8_1};
  assign _zz_biasInTemp_8_3 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_2 = {{8{_zz_biasInTemp_8_3[0]}}, _zz_biasInTemp_8_3};
  assign _zz_biasInTemp_8_5 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_4 = {{9{_zz_biasInTemp_8_5[0]}}, _zz_biasInTemp_8_5};
  assign _zz_biasInTemp_8_7 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_6 = {{10{_zz_biasInTemp_8_7[0]}}, _zz_biasInTemp_8_7};
  assign _zz_biasInTemp_8_9 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_8 = {{11{_zz_biasInTemp_8_9[0]}}, _zz_biasInTemp_8_9};
  assign _zz_biasInTemp_8_11 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_10 = {{12{_zz_biasInTemp_8_11[0]}}, _zz_biasInTemp_8_11};
  assign _zz_biasInTemp_8_13 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_12 = {{13{_zz_biasInTemp_8_13[0]}}, _zz_biasInTemp_8_13};
  assign _zz_biasInTemp_8_15 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_14 = {{14{_zz_biasInTemp_8_15[0]}}, _zz_biasInTemp_8_15};
  assign _zz_biasInTemp_8_17 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_16 = {{15{_zz_biasInTemp_8_17[0]}}, _zz_biasInTemp_8_17};
  assign _zz_biasInTemp_8_19 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_18 = {{16{_zz_biasInTemp_8_19[0]}}, _zz_biasInTemp_8_19};
  assign _zz_biasInTemp_8_21 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_20 = {{17{_zz_biasInTemp_8_21[0]}}, _zz_biasInTemp_8_21};
  assign _zz_biasInTemp_8_23 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_22 = {{18{_zz_biasInTemp_8_23[0]}}, _zz_biasInTemp_8_23};
  assign _zz_biasInTemp_8_25 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_24 = {{19{_zz_biasInTemp_8_25[0]}}, _zz_biasInTemp_8_25};
  assign _zz_biasInTemp_8_27 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_26 = {{20{_zz_biasInTemp_8_27[0]}}, _zz_biasInTemp_8_27};
  assign _zz_biasInTemp_8_29 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_28 = {{21{_zz_biasInTemp_8_29[0]}}, _zz_biasInTemp_8_29};
  assign _zz_biasInTemp_8_31 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_30 = {{22{_zz_biasInTemp_8_31[0]}}, _zz_biasInTemp_8_31};
  assign _zz_biasInTemp_8_33 = Bias_quan_8[31];
  assign _zz_biasInTemp_8_32 = {{23{_zz_biasInTemp_8_33[0]}}, _zz_biasInTemp_8_33};
  assign _zz_dataInTemp_9 = 16'h0;
  assign _zz_biasInTemp_9_1 = Bias_quan_9[31];
  assign _zz_biasInTemp_9 = {{7{_zz_biasInTemp_9_1[0]}}, _zz_biasInTemp_9_1};
  assign _zz_biasInTemp_9_3 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_2 = {{8{_zz_biasInTemp_9_3[0]}}, _zz_biasInTemp_9_3};
  assign _zz_biasInTemp_9_5 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_4 = {{9{_zz_biasInTemp_9_5[0]}}, _zz_biasInTemp_9_5};
  assign _zz_biasInTemp_9_7 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_6 = {{10{_zz_biasInTemp_9_7[0]}}, _zz_biasInTemp_9_7};
  assign _zz_biasInTemp_9_9 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_8 = {{11{_zz_biasInTemp_9_9[0]}}, _zz_biasInTemp_9_9};
  assign _zz_biasInTemp_9_11 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_10 = {{12{_zz_biasInTemp_9_11[0]}}, _zz_biasInTemp_9_11};
  assign _zz_biasInTemp_9_13 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_12 = {{13{_zz_biasInTemp_9_13[0]}}, _zz_biasInTemp_9_13};
  assign _zz_biasInTemp_9_15 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_14 = {{14{_zz_biasInTemp_9_15[0]}}, _zz_biasInTemp_9_15};
  assign _zz_biasInTemp_9_17 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_16 = {{15{_zz_biasInTemp_9_17[0]}}, _zz_biasInTemp_9_17};
  assign _zz_biasInTemp_9_19 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_18 = {{16{_zz_biasInTemp_9_19[0]}}, _zz_biasInTemp_9_19};
  assign _zz_biasInTemp_9_21 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_20 = {{17{_zz_biasInTemp_9_21[0]}}, _zz_biasInTemp_9_21};
  assign _zz_biasInTemp_9_23 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_22 = {{18{_zz_biasInTemp_9_23[0]}}, _zz_biasInTemp_9_23};
  assign _zz_biasInTemp_9_25 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_24 = {{19{_zz_biasInTemp_9_25[0]}}, _zz_biasInTemp_9_25};
  assign _zz_biasInTemp_9_27 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_26 = {{20{_zz_biasInTemp_9_27[0]}}, _zz_biasInTemp_9_27};
  assign _zz_biasInTemp_9_29 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_28 = {{21{_zz_biasInTemp_9_29[0]}}, _zz_biasInTemp_9_29};
  assign _zz_biasInTemp_9_31 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_30 = {{22{_zz_biasInTemp_9_31[0]}}, _zz_biasInTemp_9_31};
  assign _zz_biasInTemp_9_33 = Bias_quan_9[31];
  assign _zz_biasInTemp_9_32 = {{23{_zz_biasInTemp_9_33[0]}}, _zz_biasInTemp_9_33};
  assign _zz_dataInTemp_10 = 16'h0;
  assign _zz_biasInTemp_10_1 = Bias_quan_10[31];
  assign _zz_biasInTemp_10 = {{7{_zz_biasInTemp_10_1[0]}}, _zz_biasInTemp_10_1};
  assign _zz_biasInTemp_10_3 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_2 = {{8{_zz_biasInTemp_10_3[0]}}, _zz_biasInTemp_10_3};
  assign _zz_biasInTemp_10_5 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_4 = {{9{_zz_biasInTemp_10_5[0]}}, _zz_biasInTemp_10_5};
  assign _zz_biasInTemp_10_7 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_6 = {{10{_zz_biasInTemp_10_7[0]}}, _zz_biasInTemp_10_7};
  assign _zz_biasInTemp_10_9 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_8 = {{11{_zz_biasInTemp_10_9[0]}}, _zz_biasInTemp_10_9};
  assign _zz_biasInTemp_10_11 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_10 = {{12{_zz_biasInTemp_10_11[0]}}, _zz_biasInTemp_10_11};
  assign _zz_biasInTemp_10_13 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_12 = {{13{_zz_biasInTemp_10_13[0]}}, _zz_biasInTemp_10_13};
  assign _zz_biasInTemp_10_15 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_14 = {{14{_zz_biasInTemp_10_15[0]}}, _zz_biasInTemp_10_15};
  assign _zz_biasInTemp_10_17 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_16 = {{15{_zz_biasInTemp_10_17[0]}}, _zz_biasInTemp_10_17};
  assign _zz_biasInTemp_10_19 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_18 = {{16{_zz_biasInTemp_10_19[0]}}, _zz_biasInTemp_10_19};
  assign _zz_biasInTemp_10_21 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_20 = {{17{_zz_biasInTemp_10_21[0]}}, _zz_biasInTemp_10_21};
  assign _zz_biasInTemp_10_23 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_22 = {{18{_zz_biasInTemp_10_23[0]}}, _zz_biasInTemp_10_23};
  assign _zz_biasInTemp_10_25 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_24 = {{19{_zz_biasInTemp_10_25[0]}}, _zz_biasInTemp_10_25};
  assign _zz_biasInTemp_10_27 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_26 = {{20{_zz_biasInTemp_10_27[0]}}, _zz_biasInTemp_10_27};
  assign _zz_biasInTemp_10_29 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_28 = {{21{_zz_biasInTemp_10_29[0]}}, _zz_biasInTemp_10_29};
  assign _zz_biasInTemp_10_31 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_30 = {{22{_zz_biasInTemp_10_31[0]}}, _zz_biasInTemp_10_31};
  assign _zz_biasInTemp_10_33 = Bias_quan_10[31];
  assign _zz_biasInTemp_10_32 = {{23{_zz_biasInTemp_10_33[0]}}, _zz_biasInTemp_10_33};
  assign _zz_dataInTemp_11 = 16'h0;
  assign _zz_biasInTemp_11_1 = Bias_quan_11[31];
  assign _zz_biasInTemp_11 = {{7{_zz_biasInTemp_11_1[0]}}, _zz_biasInTemp_11_1};
  assign _zz_biasInTemp_11_3 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_2 = {{8{_zz_biasInTemp_11_3[0]}}, _zz_biasInTemp_11_3};
  assign _zz_biasInTemp_11_5 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_4 = {{9{_zz_biasInTemp_11_5[0]}}, _zz_biasInTemp_11_5};
  assign _zz_biasInTemp_11_7 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_6 = {{10{_zz_biasInTemp_11_7[0]}}, _zz_biasInTemp_11_7};
  assign _zz_biasInTemp_11_9 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_8 = {{11{_zz_biasInTemp_11_9[0]}}, _zz_biasInTemp_11_9};
  assign _zz_biasInTemp_11_11 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_10 = {{12{_zz_biasInTemp_11_11[0]}}, _zz_biasInTemp_11_11};
  assign _zz_biasInTemp_11_13 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_12 = {{13{_zz_biasInTemp_11_13[0]}}, _zz_biasInTemp_11_13};
  assign _zz_biasInTemp_11_15 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_14 = {{14{_zz_biasInTemp_11_15[0]}}, _zz_biasInTemp_11_15};
  assign _zz_biasInTemp_11_17 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_16 = {{15{_zz_biasInTemp_11_17[0]}}, _zz_biasInTemp_11_17};
  assign _zz_biasInTemp_11_19 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_18 = {{16{_zz_biasInTemp_11_19[0]}}, _zz_biasInTemp_11_19};
  assign _zz_biasInTemp_11_21 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_20 = {{17{_zz_biasInTemp_11_21[0]}}, _zz_biasInTemp_11_21};
  assign _zz_biasInTemp_11_23 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_22 = {{18{_zz_biasInTemp_11_23[0]}}, _zz_biasInTemp_11_23};
  assign _zz_biasInTemp_11_25 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_24 = {{19{_zz_biasInTemp_11_25[0]}}, _zz_biasInTemp_11_25};
  assign _zz_biasInTemp_11_27 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_26 = {{20{_zz_biasInTemp_11_27[0]}}, _zz_biasInTemp_11_27};
  assign _zz_biasInTemp_11_29 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_28 = {{21{_zz_biasInTemp_11_29[0]}}, _zz_biasInTemp_11_29};
  assign _zz_biasInTemp_11_31 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_30 = {{22{_zz_biasInTemp_11_31[0]}}, _zz_biasInTemp_11_31};
  assign _zz_biasInTemp_11_33 = Bias_quan_11[31];
  assign _zz_biasInTemp_11_32 = {{23{_zz_biasInTemp_11_33[0]}}, _zz_biasInTemp_11_33};
  assign _zz_dataInTemp_12 = 16'h0;
  assign _zz_biasInTemp_12_1 = Bias_quan_12[31];
  assign _zz_biasInTemp_12 = {{7{_zz_biasInTemp_12_1[0]}}, _zz_biasInTemp_12_1};
  assign _zz_biasInTemp_12_3 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_2 = {{8{_zz_biasInTemp_12_3[0]}}, _zz_biasInTemp_12_3};
  assign _zz_biasInTemp_12_5 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_4 = {{9{_zz_biasInTemp_12_5[0]}}, _zz_biasInTemp_12_5};
  assign _zz_biasInTemp_12_7 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_6 = {{10{_zz_biasInTemp_12_7[0]}}, _zz_biasInTemp_12_7};
  assign _zz_biasInTemp_12_9 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_8 = {{11{_zz_biasInTemp_12_9[0]}}, _zz_biasInTemp_12_9};
  assign _zz_biasInTemp_12_11 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_10 = {{12{_zz_biasInTemp_12_11[0]}}, _zz_biasInTemp_12_11};
  assign _zz_biasInTemp_12_13 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_12 = {{13{_zz_biasInTemp_12_13[0]}}, _zz_biasInTemp_12_13};
  assign _zz_biasInTemp_12_15 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_14 = {{14{_zz_biasInTemp_12_15[0]}}, _zz_biasInTemp_12_15};
  assign _zz_biasInTemp_12_17 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_16 = {{15{_zz_biasInTemp_12_17[0]}}, _zz_biasInTemp_12_17};
  assign _zz_biasInTemp_12_19 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_18 = {{16{_zz_biasInTemp_12_19[0]}}, _zz_biasInTemp_12_19};
  assign _zz_biasInTemp_12_21 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_20 = {{17{_zz_biasInTemp_12_21[0]}}, _zz_biasInTemp_12_21};
  assign _zz_biasInTemp_12_23 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_22 = {{18{_zz_biasInTemp_12_23[0]}}, _zz_biasInTemp_12_23};
  assign _zz_biasInTemp_12_25 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_24 = {{19{_zz_biasInTemp_12_25[0]}}, _zz_biasInTemp_12_25};
  assign _zz_biasInTemp_12_27 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_26 = {{20{_zz_biasInTemp_12_27[0]}}, _zz_biasInTemp_12_27};
  assign _zz_biasInTemp_12_29 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_28 = {{21{_zz_biasInTemp_12_29[0]}}, _zz_biasInTemp_12_29};
  assign _zz_biasInTemp_12_31 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_30 = {{22{_zz_biasInTemp_12_31[0]}}, _zz_biasInTemp_12_31};
  assign _zz_biasInTemp_12_33 = Bias_quan_12[31];
  assign _zz_biasInTemp_12_32 = {{23{_zz_biasInTemp_12_33[0]}}, _zz_biasInTemp_12_33};
  assign _zz_dataInTemp_13 = 16'h0;
  assign _zz_biasInTemp_13_1 = Bias_quan_13[31];
  assign _zz_biasInTemp_13 = {{7{_zz_biasInTemp_13_1[0]}}, _zz_biasInTemp_13_1};
  assign _zz_biasInTemp_13_3 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_2 = {{8{_zz_biasInTemp_13_3[0]}}, _zz_biasInTemp_13_3};
  assign _zz_biasInTemp_13_5 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_4 = {{9{_zz_biasInTemp_13_5[0]}}, _zz_biasInTemp_13_5};
  assign _zz_biasInTemp_13_7 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_6 = {{10{_zz_biasInTemp_13_7[0]}}, _zz_biasInTemp_13_7};
  assign _zz_biasInTemp_13_9 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_8 = {{11{_zz_biasInTemp_13_9[0]}}, _zz_biasInTemp_13_9};
  assign _zz_biasInTemp_13_11 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_10 = {{12{_zz_biasInTemp_13_11[0]}}, _zz_biasInTemp_13_11};
  assign _zz_biasInTemp_13_13 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_12 = {{13{_zz_biasInTemp_13_13[0]}}, _zz_biasInTemp_13_13};
  assign _zz_biasInTemp_13_15 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_14 = {{14{_zz_biasInTemp_13_15[0]}}, _zz_biasInTemp_13_15};
  assign _zz_biasInTemp_13_17 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_16 = {{15{_zz_biasInTemp_13_17[0]}}, _zz_biasInTemp_13_17};
  assign _zz_biasInTemp_13_19 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_18 = {{16{_zz_biasInTemp_13_19[0]}}, _zz_biasInTemp_13_19};
  assign _zz_biasInTemp_13_21 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_20 = {{17{_zz_biasInTemp_13_21[0]}}, _zz_biasInTemp_13_21};
  assign _zz_biasInTemp_13_23 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_22 = {{18{_zz_biasInTemp_13_23[0]}}, _zz_biasInTemp_13_23};
  assign _zz_biasInTemp_13_25 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_24 = {{19{_zz_biasInTemp_13_25[0]}}, _zz_biasInTemp_13_25};
  assign _zz_biasInTemp_13_27 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_26 = {{20{_zz_biasInTemp_13_27[0]}}, _zz_biasInTemp_13_27};
  assign _zz_biasInTemp_13_29 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_28 = {{21{_zz_biasInTemp_13_29[0]}}, _zz_biasInTemp_13_29};
  assign _zz_biasInTemp_13_31 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_30 = {{22{_zz_biasInTemp_13_31[0]}}, _zz_biasInTemp_13_31};
  assign _zz_biasInTemp_13_33 = Bias_quan_13[31];
  assign _zz_biasInTemp_13_32 = {{23{_zz_biasInTemp_13_33[0]}}, _zz_biasInTemp_13_33};
  assign _zz_dataInTemp_14 = 16'h0;
  assign _zz_biasInTemp_14_1 = Bias_quan_14[31];
  assign _zz_biasInTemp_14 = {{7{_zz_biasInTemp_14_1[0]}}, _zz_biasInTemp_14_1};
  assign _zz_biasInTemp_14_3 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_2 = {{8{_zz_biasInTemp_14_3[0]}}, _zz_biasInTemp_14_3};
  assign _zz_biasInTemp_14_5 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_4 = {{9{_zz_biasInTemp_14_5[0]}}, _zz_biasInTemp_14_5};
  assign _zz_biasInTemp_14_7 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_6 = {{10{_zz_biasInTemp_14_7[0]}}, _zz_biasInTemp_14_7};
  assign _zz_biasInTemp_14_9 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_8 = {{11{_zz_biasInTemp_14_9[0]}}, _zz_biasInTemp_14_9};
  assign _zz_biasInTemp_14_11 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_10 = {{12{_zz_biasInTemp_14_11[0]}}, _zz_biasInTemp_14_11};
  assign _zz_biasInTemp_14_13 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_12 = {{13{_zz_biasInTemp_14_13[0]}}, _zz_biasInTemp_14_13};
  assign _zz_biasInTemp_14_15 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_14 = {{14{_zz_biasInTemp_14_15[0]}}, _zz_biasInTemp_14_15};
  assign _zz_biasInTemp_14_17 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_16 = {{15{_zz_biasInTemp_14_17[0]}}, _zz_biasInTemp_14_17};
  assign _zz_biasInTemp_14_19 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_18 = {{16{_zz_biasInTemp_14_19[0]}}, _zz_biasInTemp_14_19};
  assign _zz_biasInTemp_14_21 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_20 = {{17{_zz_biasInTemp_14_21[0]}}, _zz_biasInTemp_14_21};
  assign _zz_biasInTemp_14_23 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_22 = {{18{_zz_biasInTemp_14_23[0]}}, _zz_biasInTemp_14_23};
  assign _zz_biasInTemp_14_25 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_24 = {{19{_zz_biasInTemp_14_25[0]}}, _zz_biasInTemp_14_25};
  assign _zz_biasInTemp_14_27 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_26 = {{20{_zz_biasInTemp_14_27[0]}}, _zz_biasInTemp_14_27};
  assign _zz_biasInTemp_14_29 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_28 = {{21{_zz_biasInTemp_14_29[0]}}, _zz_biasInTemp_14_29};
  assign _zz_biasInTemp_14_31 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_30 = {{22{_zz_biasInTemp_14_31[0]}}, _zz_biasInTemp_14_31};
  assign _zz_biasInTemp_14_33 = Bias_quan_14[31];
  assign _zz_biasInTemp_14_32 = {{23{_zz_biasInTemp_14_33[0]}}, _zz_biasInTemp_14_33};
  assign _zz_dataInTemp_15 = 16'h0;
  assign _zz_biasInTemp_15_1 = Bias_quan_15[31];
  assign _zz_biasInTemp_15 = {{7{_zz_biasInTemp_15_1[0]}}, _zz_biasInTemp_15_1};
  assign _zz_biasInTemp_15_3 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_2 = {{8{_zz_biasInTemp_15_3[0]}}, _zz_biasInTemp_15_3};
  assign _zz_biasInTemp_15_5 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_4 = {{9{_zz_biasInTemp_15_5[0]}}, _zz_biasInTemp_15_5};
  assign _zz_biasInTemp_15_7 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_6 = {{10{_zz_biasInTemp_15_7[0]}}, _zz_biasInTemp_15_7};
  assign _zz_biasInTemp_15_9 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_8 = {{11{_zz_biasInTemp_15_9[0]}}, _zz_biasInTemp_15_9};
  assign _zz_biasInTemp_15_11 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_10 = {{12{_zz_biasInTemp_15_11[0]}}, _zz_biasInTemp_15_11};
  assign _zz_biasInTemp_15_13 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_12 = {{13{_zz_biasInTemp_15_13[0]}}, _zz_biasInTemp_15_13};
  assign _zz_biasInTemp_15_15 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_14 = {{14{_zz_biasInTemp_15_15[0]}}, _zz_biasInTemp_15_15};
  assign _zz_biasInTemp_15_17 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_16 = {{15{_zz_biasInTemp_15_17[0]}}, _zz_biasInTemp_15_17};
  assign _zz_biasInTemp_15_19 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_18 = {{16{_zz_biasInTemp_15_19[0]}}, _zz_biasInTemp_15_19};
  assign _zz_biasInTemp_15_21 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_20 = {{17{_zz_biasInTemp_15_21[0]}}, _zz_biasInTemp_15_21};
  assign _zz_biasInTemp_15_23 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_22 = {{18{_zz_biasInTemp_15_23[0]}}, _zz_biasInTemp_15_23};
  assign _zz_biasInTemp_15_25 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_24 = {{19{_zz_biasInTemp_15_25[0]}}, _zz_biasInTemp_15_25};
  assign _zz_biasInTemp_15_27 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_26 = {{20{_zz_biasInTemp_15_27[0]}}, _zz_biasInTemp_15_27};
  assign _zz_biasInTemp_15_29 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_28 = {{21{_zz_biasInTemp_15_29[0]}}, _zz_biasInTemp_15_29};
  assign _zz_biasInTemp_15_31 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_30 = {{22{_zz_biasInTemp_15_31[0]}}, _zz_biasInTemp_15_31};
  assign _zz_biasInTemp_15_33 = Bias_quan_15[31];
  assign _zz_biasInTemp_15_32 = {{23{_zz_biasInTemp_15_33[0]}}, _zz_biasInTemp_15_33};
  biasAdd addSub (
    .A   (dataInTemp_0[47:0]), //i
    .B   (biasInTemp_0[47:0]), //i
    .S   (addSub_S[47:0]    ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_1 (
    .A   (dataInTemp_1[47:0]), //i
    .B   (biasInTemp_1[47:0]), //i
    .S   (addSub_1_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_2 (
    .A   (dataInTemp_2[47:0]), //i
    .B   (biasInTemp_2[47:0]), //i
    .S   (addSub_2_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_3 (
    .A   (dataInTemp_3[47:0]), //i
    .B   (biasInTemp_3[47:0]), //i
    .S   (addSub_3_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_4 (
    .A   (dataInTemp_4[47:0]), //i
    .B   (biasInTemp_4[47:0]), //i
    .S   (addSub_4_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_5 (
    .A   (dataInTemp_5[47:0]), //i
    .B   (biasInTemp_5[47:0]), //i
    .S   (addSub_5_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_6 (
    .A   (dataInTemp_6[47:0]), //i
    .B   (biasInTemp_6[47:0]), //i
    .S   (addSub_6_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_7 (
    .A   (dataInTemp_7[47:0]), //i
    .B   (biasInTemp_7[47:0]), //i
    .S   (addSub_7_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_8 (
    .A   (dataInTemp_8[47:0]), //i
    .B   (biasInTemp_8[47:0]), //i
    .S   (addSub_8_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_9 (
    .A   (dataInTemp_9[47:0]), //i
    .B   (biasInTemp_9[47:0]), //i
    .S   (addSub_9_S[47:0]  ), //o
    .CLK (clk               )  //i
  );
  biasAdd addSub_10 (
    .A   (dataInTemp_10[47:0]), //i
    .B   (biasInTemp_10[47:0]), //i
    .S   (addSub_10_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  biasAdd addSub_11 (
    .A   (dataInTemp_11[47:0]), //i
    .B   (biasInTemp_11[47:0]), //i
    .S   (addSub_11_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  biasAdd addSub_12 (
    .A   (dataInTemp_12[47:0]), //i
    .B   (biasInTemp_12[47:0]), //i
    .S   (addSub_12_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  biasAdd addSub_13 (
    .A   (dataInTemp_13[47:0]), //i
    .B   (biasInTemp_13[47:0]), //i
    .S   (addSub_13_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  biasAdd addSub_14 (
    .A   (dataInTemp_14[47:0]), //i
    .B   (biasInTemp_14[47:0]), //i
    .S   (addSub_14_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  biasAdd addSub_15 (
    .A   (dataInTemp_15[47:0]), //i
    .B   (biasInTemp_15[47:0]), //i
    .S   (addSub_15_S[47:0]  ), //o
    .CLK (clk                )  //i
  );
  assign switch_Quan_l67 = Bias_quan_0[30 : 24];
  assign switch_Quan_l67_1 = Bias_quan_1[30 : 24];
  assign switch_Quan_l67_2 = Bias_quan_2[30 : 24];
  assign switch_Quan_l67_3 = Bias_quan_3[30 : 24];
  assign switch_Quan_l67_4 = Bias_quan_4[30 : 24];
  assign switch_Quan_l67_5 = Bias_quan_5[30 : 24];
  assign switch_Quan_l67_6 = Bias_quan_6[30 : 24];
  assign switch_Quan_l67_7 = Bias_quan_7[30 : 24];
  assign switch_Quan_l67_8 = Bias_quan_8[30 : 24];
  assign switch_Quan_l67_9 = Bias_quan_9[30 : 24];
  assign switch_Quan_l67_10 = Bias_quan_10[30 : 24];
  assign switch_Quan_l67_11 = Bias_quan_11[30 : 24];
  assign switch_Quan_l67_12 = Bias_quan_12[30 : 24];
  assign switch_Quan_l67_13 = Bias_quan_13[30 : 24];
  assign switch_Quan_l67_14 = Bias_quan_14[30 : 24];
  assign switch_Quan_l67_15 = Bias_quan_15[30 : 24];
  assign Bias_dataOut_0 = addSub_S;
  assign Bias_dataOut_1 = addSub_1_S;
  assign Bias_dataOut_2 = addSub_2_S;
  assign Bias_dataOut_3 = addSub_3_S;
  assign Bias_dataOut_4 = addSub_4_S;
  assign Bias_dataOut_5 = addSub_5_S;
  assign Bias_dataOut_6 = addSub_6_S;
  assign Bias_dataOut_7 = addSub_7_S;
  assign Bias_dataOut_8 = addSub_8_S;
  assign Bias_dataOut_9 = addSub_9_S;
  assign Bias_dataOut_10 = addSub_10_S;
  assign Bias_dataOut_11 = addSub_11_S;
  assign Bias_dataOut_12 = addSub_12_S;
  assign Bias_dataOut_13 = addSub_13_S;
  assign Bias_dataOut_14 = addSub_14_S;
  assign Bias_dataOut_15 = addSub_15_S;
  always @(posedge clk) begin
    dataInTemp_0 <= {Bias_dataIn_0,_zz_dataInTemp_0};
    case(switch_Quan_l67)
      7'h0 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0,Bias_quan_0[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_2,Bias_quan_0[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_4,Bias_quan_0[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_6,Bias_quan_0[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_8,Bias_quan_0[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_10,Bias_quan_0[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_12,Bias_quan_0[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_14,Bias_quan_0[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_16,Bias_quan_0[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_18,Bias_quan_0[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_20,Bias_quan_0[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_22,Bias_quan_0[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_24,Bias_quan_0[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_26,Bias_quan_0[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_28,Bias_quan_0[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_0 <= {{_zz_biasInTemp_0_30,Bias_quan_0[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_0 <= {_zz_biasInTemp_0_32,Bias_quan_0[23 : 0]};
      end
      default : begin
        biasInTemp_0 <= 48'h0;
      end
    endcase
    dataInTemp_1 <= {Bias_dataIn_1,_zz_dataInTemp_1};
    case(switch_Quan_l67_1)
      7'h0 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1,Bias_quan_1[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_2,Bias_quan_1[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_4,Bias_quan_1[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_6,Bias_quan_1[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_8,Bias_quan_1[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_10,Bias_quan_1[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_12,Bias_quan_1[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_14,Bias_quan_1[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_16,Bias_quan_1[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_18,Bias_quan_1[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_20,Bias_quan_1[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_22,Bias_quan_1[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_24,Bias_quan_1[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_26,Bias_quan_1[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_28,Bias_quan_1[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_1 <= {{_zz_biasInTemp_1_30,Bias_quan_1[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_1 <= {_zz_biasInTemp_1_32,Bias_quan_1[23 : 0]};
      end
      default : begin
        biasInTemp_1 <= 48'h0;
      end
    endcase
    dataInTemp_2 <= {Bias_dataIn_2,_zz_dataInTemp_2};
    case(switch_Quan_l67_2)
      7'h0 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2,Bias_quan_2[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_2,Bias_quan_2[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_4,Bias_quan_2[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_6,Bias_quan_2[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_8,Bias_quan_2[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_10,Bias_quan_2[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_12,Bias_quan_2[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_14,Bias_quan_2[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_16,Bias_quan_2[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_18,Bias_quan_2[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_20,Bias_quan_2[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_22,Bias_quan_2[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_24,Bias_quan_2[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_26,Bias_quan_2[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_28,Bias_quan_2[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_2 <= {{_zz_biasInTemp_2_30,Bias_quan_2[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_2 <= {_zz_biasInTemp_2_32,Bias_quan_2[23 : 0]};
      end
      default : begin
        biasInTemp_2 <= 48'h0;
      end
    endcase
    dataInTemp_3 <= {Bias_dataIn_3,_zz_dataInTemp_3};
    case(switch_Quan_l67_3)
      7'h0 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3,Bias_quan_3[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_2,Bias_quan_3[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_4,Bias_quan_3[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_6,Bias_quan_3[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_8,Bias_quan_3[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_10,Bias_quan_3[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_12,Bias_quan_3[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_14,Bias_quan_3[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_16,Bias_quan_3[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_18,Bias_quan_3[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_20,Bias_quan_3[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_22,Bias_quan_3[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_24,Bias_quan_3[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_26,Bias_quan_3[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_28,Bias_quan_3[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_3 <= {{_zz_biasInTemp_3_30,Bias_quan_3[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_3 <= {_zz_biasInTemp_3_32,Bias_quan_3[23 : 0]};
      end
      default : begin
        biasInTemp_3 <= 48'h0;
      end
    endcase
    dataInTemp_4 <= {Bias_dataIn_4,_zz_dataInTemp_4};
    case(switch_Quan_l67_4)
      7'h0 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4,Bias_quan_4[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_2,Bias_quan_4[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_4,Bias_quan_4[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_6,Bias_quan_4[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_8,Bias_quan_4[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_10,Bias_quan_4[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_12,Bias_quan_4[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_14,Bias_quan_4[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_16,Bias_quan_4[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_18,Bias_quan_4[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_20,Bias_quan_4[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_22,Bias_quan_4[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_24,Bias_quan_4[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_26,Bias_quan_4[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_28,Bias_quan_4[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_4 <= {{_zz_biasInTemp_4_30,Bias_quan_4[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_4 <= {_zz_biasInTemp_4_32,Bias_quan_4[23 : 0]};
      end
      default : begin
        biasInTemp_4 <= 48'h0;
      end
    endcase
    dataInTemp_5 <= {Bias_dataIn_5,_zz_dataInTemp_5};
    case(switch_Quan_l67_5)
      7'h0 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5,Bias_quan_5[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_2,Bias_quan_5[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_4,Bias_quan_5[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_6,Bias_quan_5[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_8,Bias_quan_5[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_10,Bias_quan_5[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_12,Bias_quan_5[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_14,Bias_quan_5[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_16,Bias_quan_5[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_18,Bias_quan_5[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_20,Bias_quan_5[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_22,Bias_quan_5[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_24,Bias_quan_5[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_26,Bias_quan_5[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_28,Bias_quan_5[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_5 <= {{_zz_biasInTemp_5_30,Bias_quan_5[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_5 <= {_zz_biasInTemp_5_32,Bias_quan_5[23 : 0]};
      end
      default : begin
        biasInTemp_5 <= 48'h0;
      end
    endcase
    dataInTemp_6 <= {Bias_dataIn_6,_zz_dataInTemp_6};
    case(switch_Quan_l67_6)
      7'h0 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6,Bias_quan_6[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_2,Bias_quan_6[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_4,Bias_quan_6[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_6,Bias_quan_6[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_8,Bias_quan_6[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_10,Bias_quan_6[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_12,Bias_quan_6[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_14,Bias_quan_6[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_16,Bias_quan_6[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_18,Bias_quan_6[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_20,Bias_quan_6[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_22,Bias_quan_6[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_24,Bias_quan_6[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_26,Bias_quan_6[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_28,Bias_quan_6[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_6 <= {{_zz_biasInTemp_6_30,Bias_quan_6[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_6 <= {_zz_biasInTemp_6_32,Bias_quan_6[23 : 0]};
      end
      default : begin
        biasInTemp_6 <= 48'h0;
      end
    endcase
    dataInTemp_7 <= {Bias_dataIn_7,_zz_dataInTemp_7};
    case(switch_Quan_l67_7)
      7'h0 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7,Bias_quan_7[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_2,Bias_quan_7[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_4,Bias_quan_7[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_6,Bias_quan_7[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_8,Bias_quan_7[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_10,Bias_quan_7[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_12,Bias_quan_7[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_14,Bias_quan_7[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_16,Bias_quan_7[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_18,Bias_quan_7[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_20,Bias_quan_7[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_22,Bias_quan_7[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_24,Bias_quan_7[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_26,Bias_quan_7[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_28,Bias_quan_7[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_7 <= {{_zz_biasInTemp_7_30,Bias_quan_7[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_7 <= {_zz_biasInTemp_7_32,Bias_quan_7[23 : 0]};
      end
      default : begin
        biasInTemp_7 <= 48'h0;
      end
    endcase
    dataInTemp_8 <= {Bias_dataIn_8,_zz_dataInTemp_8};
    case(switch_Quan_l67_8)
      7'h0 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8,Bias_quan_8[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_2,Bias_quan_8[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_4,Bias_quan_8[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_6,Bias_quan_8[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_8,Bias_quan_8[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_10,Bias_quan_8[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_12,Bias_quan_8[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_14,Bias_quan_8[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_16,Bias_quan_8[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_18,Bias_quan_8[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_20,Bias_quan_8[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_22,Bias_quan_8[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_24,Bias_quan_8[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_26,Bias_quan_8[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_28,Bias_quan_8[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_8 <= {{_zz_biasInTemp_8_30,Bias_quan_8[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_8 <= {_zz_biasInTemp_8_32,Bias_quan_8[23 : 0]};
      end
      default : begin
        biasInTemp_8 <= 48'h0;
      end
    endcase
    dataInTemp_9 <= {Bias_dataIn_9,_zz_dataInTemp_9};
    case(switch_Quan_l67_9)
      7'h0 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9,Bias_quan_9[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_2,Bias_quan_9[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_4,Bias_quan_9[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_6,Bias_quan_9[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_8,Bias_quan_9[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_10,Bias_quan_9[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_12,Bias_quan_9[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_14,Bias_quan_9[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_16,Bias_quan_9[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_18,Bias_quan_9[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_20,Bias_quan_9[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_22,Bias_quan_9[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_24,Bias_quan_9[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_26,Bias_quan_9[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_28,Bias_quan_9[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_9 <= {{_zz_biasInTemp_9_30,Bias_quan_9[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_9 <= {_zz_biasInTemp_9_32,Bias_quan_9[23 : 0]};
      end
      default : begin
        biasInTemp_9 <= 48'h0;
      end
    endcase
    dataInTemp_10 <= {Bias_dataIn_10,_zz_dataInTemp_10};
    case(switch_Quan_l67_10)
      7'h0 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10,Bias_quan_10[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_2,Bias_quan_10[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_4,Bias_quan_10[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_6,Bias_quan_10[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_8,Bias_quan_10[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_10,Bias_quan_10[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_12,Bias_quan_10[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_14,Bias_quan_10[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_16,Bias_quan_10[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_18,Bias_quan_10[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_20,Bias_quan_10[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_22,Bias_quan_10[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_24,Bias_quan_10[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_26,Bias_quan_10[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_28,Bias_quan_10[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_10 <= {{_zz_biasInTemp_10_30,Bias_quan_10[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_10 <= {_zz_biasInTemp_10_32,Bias_quan_10[23 : 0]};
      end
      default : begin
        biasInTemp_10 <= 48'h0;
      end
    endcase
    dataInTemp_11 <= {Bias_dataIn_11,_zz_dataInTemp_11};
    case(switch_Quan_l67_11)
      7'h0 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11,Bias_quan_11[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_2,Bias_quan_11[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_4,Bias_quan_11[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_6,Bias_quan_11[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_8,Bias_quan_11[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_10,Bias_quan_11[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_12,Bias_quan_11[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_14,Bias_quan_11[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_16,Bias_quan_11[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_18,Bias_quan_11[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_20,Bias_quan_11[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_22,Bias_quan_11[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_24,Bias_quan_11[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_26,Bias_quan_11[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_28,Bias_quan_11[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_11 <= {{_zz_biasInTemp_11_30,Bias_quan_11[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_11 <= {_zz_biasInTemp_11_32,Bias_quan_11[23 : 0]};
      end
      default : begin
        biasInTemp_11 <= 48'h0;
      end
    endcase
    dataInTemp_12 <= {Bias_dataIn_12,_zz_dataInTemp_12};
    case(switch_Quan_l67_12)
      7'h0 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12,Bias_quan_12[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_2,Bias_quan_12[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_4,Bias_quan_12[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_6,Bias_quan_12[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_8,Bias_quan_12[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_10,Bias_quan_12[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_12,Bias_quan_12[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_14,Bias_quan_12[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_16,Bias_quan_12[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_18,Bias_quan_12[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_20,Bias_quan_12[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_22,Bias_quan_12[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_24,Bias_quan_12[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_26,Bias_quan_12[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_28,Bias_quan_12[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_12 <= {{_zz_biasInTemp_12_30,Bias_quan_12[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_12 <= {_zz_biasInTemp_12_32,Bias_quan_12[23 : 0]};
      end
      default : begin
        biasInTemp_12 <= 48'h0;
      end
    endcase
    dataInTemp_13 <= {Bias_dataIn_13,_zz_dataInTemp_13};
    case(switch_Quan_l67_13)
      7'h0 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13,Bias_quan_13[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_2,Bias_quan_13[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_4,Bias_quan_13[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_6,Bias_quan_13[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_8,Bias_quan_13[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_10,Bias_quan_13[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_12,Bias_quan_13[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_14,Bias_quan_13[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_16,Bias_quan_13[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_18,Bias_quan_13[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_20,Bias_quan_13[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_22,Bias_quan_13[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_24,Bias_quan_13[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_26,Bias_quan_13[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_28,Bias_quan_13[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_13 <= {{_zz_biasInTemp_13_30,Bias_quan_13[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_13 <= {_zz_biasInTemp_13_32,Bias_quan_13[23 : 0]};
      end
      default : begin
        biasInTemp_13 <= 48'h0;
      end
    endcase
    dataInTemp_14 <= {Bias_dataIn_14,_zz_dataInTemp_14};
    case(switch_Quan_l67_14)
      7'h0 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14,Bias_quan_14[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_2,Bias_quan_14[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_4,Bias_quan_14[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_6,Bias_quan_14[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_8,Bias_quan_14[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_10,Bias_quan_14[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_12,Bias_quan_14[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_14,Bias_quan_14[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_16,Bias_quan_14[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_18,Bias_quan_14[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_20,Bias_quan_14[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_22,Bias_quan_14[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_24,Bias_quan_14[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_26,Bias_quan_14[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_28,Bias_quan_14[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_14 <= {{_zz_biasInTemp_14_30,Bias_quan_14[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_14 <= {_zz_biasInTemp_14_32,Bias_quan_14[23 : 0]};
      end
      default : begin
        biasInTemp_14 <= 48'h0;
      end
    endcase
    dataInTemp_15 <= {Bias_dataIn_15,_zz_dataInTemp_15};
    case(switch_Quan_l67_15)
      7'h0 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15,Bias_quan_15[23 : 0]},16'h0};
      end
      7'h01 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_2,Bias_quan_15[23 : 0]},15'h0};
      end
      7'h02 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_4,Bias_quan_15[23 : 0]},14'h0};
      end
      7'h03 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_6,Bias_quan_15[23 : 0]},13'h0};
      end
      7'h04 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_8,Bias_quan_15[23 : 0]},12'h0};
      end
      7'h05 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_10,Bias_quan_15[23 : 0]},11'h0};
      end
      7'h06 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_12,Bias_quan_15[23 : 0]},10'h0};
      end
      7'h07 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_14,Bias_quan_15[23 : 0]},9'h0};
      end
      7'h08 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_16,Bias_quan_15[23 : 0]},8'h0};
      end
      7'h09 : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_18,Bias_quan_15[23 : 0]},7'h0};
      end
      7'h0a : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_20,Bias_quan_15[23 : 0]},6'h0};
      end
      7'h0b : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_22,Bias_quan_15[23 : 0]},5'h0};
      end
      7'h0c : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_24,Bias_quan_15[23 : 0]},4'b0000};
      end
      7'h0d : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_26,Bias_quan_15[23 : 0]},3'b000};
      end
      7'h0e : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_28,Bias_quan_15[23 : 0]},2'b00};
      end
      7'h0f : begin
        biasInTemp_15 <= {{_zz_biasInTemp_15_30,Bias_quan_15[23 : 0]},1'b0};
      end
      7'h10 : begin
        biasInTemp_15 <= {_zz_biasInTemp_15_32,Bias_quan_15[23 : 0]};
      end
      default : begin
        biasInTemp_15 <= 48'h0;
      end
    endcase
  end


endmodule

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

//FifoSync_1 replaced by FifoSync_1

module FifoSync_1 (
  input               wr_en,
  input      [127:0]  din,
  output     [127:0]  dout,
  input               rd_en,
  input               reset,
  input               clk
);

  wire       [127:0]  xpm_fifo_sync_1_dout;
  wire                injectdbiterr;
  wire                injectsbiterr;
  wire                sleep;

  xpm_fifo_sync #(
    .CASCADE_HEIGHT(0),
    .DOUT_RESET_VALUE(0),
    .ECC_MODE("no_ecc"),
    .FIFO_MEMORY_TYPE("block"),
    .FIFO_READ_LATENCY(0),
    .FIFO_WRITE_DEPTH(8192),
    .FULL_RESET_VALUE(0),
    .PROG_EMPTY_THRESH(5),
    .PROG_FULL_THRESH(8187),
    .RD_DATA_COUNT_WIDTH(14),
    .READ_DATA_WIDTH(128),
    .READ_MODE("fwft"),
    .SIM_ASSERT_CHK(0),
    .USE_ADV_FEATURES("0707"),
    .WAKEUP_TIME(0),
    .WRITE_DATA_WIDTH(128),
    .WR_DATA_COUNT_WIDTH(14)
  ) xpm_fifo_sync_1 (
    .dout          (xpm_fifo_sync_1_dout[127:0]), //o
    .din           (din[127:0]                 ), //i
    .injectdbiterr (injectdbiterr              ), //i
    .injectsbiterr (injectsbiterr              ), //i
    .rd_en         (rd_en                      ), //i
    .rst           (reset                      ), //i
    .sleep         (sleep                      ), //i
    .wr_clk        (clk                        ), //i
    .wr_en         (wr_en                      )  //i
  );
  assign injectdbiterr = 1'b0;
  assign injectsbiterr = 1'b0;
  assign sleep = 1'b0;
  assign dout = xpm_fifo_sync_1_dout;

endmodule

module FifoSync (
  input               wr_en,
  input      [127:0]  din,
  output     [127:0]  dout,
  input               rd_en,
  output     [13:0]   wr_data_count,
  output     [13:0]   rd_data_count,
  input               reset,
  input               clk
);

  wire       [127:0]  xpm_fifo_sync_1_dout;
  wire       [13:0]   xpm_fifo_sync_1_rd_data_count;
  wire       [13:0]   xpm_fifo_sync_1_wr_data_count;
  wire                injectdbiterr;
  wire                injectsbiterr;
  wire                sleep;

  xpm_fifo_sync #(
    .CASCADE_HEIGHT(0),
    .DOUT_RESET_VALUE(0),
    .ECC_MODE("no_ecc"),
    .FIFO_MEMORY_TYPE("block"),
    .FIFO_READ_LATENCY(0),
    .FIFO_WRITE_DEPTH(8192),
    .FULL_RESET_VALUE(0),
    .PROG_EMPTY_THRESH(5),
    .PROG_FULL_THRESH(8187),
    .RD_DATA_COUNT_WIDTH(14),
    .READ_DATA_WIDTH(128),
    .READ_MODE("fwft"),
    .SIM_ASSERT_CHK(0),
    .USE_ADV_FEATURES("0707"),
    .WAKEUP_TIME(0),
    .WRITE_DATA_WIDTH(128),
    .WR_DATA_COUNT_WIDTH(14)
  ) xpm_fifo_sync_1 (
    .dout          (xpm_fifo_sync_1_dout[127:0]        ), //o
    .rd_data_count (xpm_fifo_sync_1_rd_data_count[13:0]), //o
    .wr_data_count (xpm_fifo_sync_1_wr_data_count[13:0]), //o
    .din           (din[127:0]                         ), //i
    .injectdbiterr (injectdbiterr                      ), //i
    .injectsbiterr (injectsbiterr                      ), //i
    .rd_en         (rd_en                              ), //i
    .rst           (reset                              ), //i
    .sleep         (sleep                              ), //i
    .wr_clk        (clk                                ), //i
    .wr_en         (wr_en                              )  //i
  );
  assign injectdbiterr = 1'b0;
  assign injectsbiterr = 1'b0;
  assign sleep = 1'b0;
  assign dout = xpm_fifo_sync_1_dout;
  assign rd_data_count = xpm_fifo_sync_1_rd_data_count;
  assign wr_data_count = xpm_fifo_sync_1_wr_data_count;

endmodule

//sdpram_144 replaced by sdpram_144

//sdpram_144 replaced by sdpram_144

module sdpram_144 (
  output     [511:0]  doutb,
  input      [7:0]    addra,
  input      [5:0]    addrb,
  input      [127:0]  dina,
  input               ena,
  input               enb,
  input      [0:0]    wea,
  input               clk
);

  wire       [511:0]  temp_doutb;
  wire                injectdbiterra;
  wire                injectsbiterra;
  wire                regceb;
  wire                rstb;
  wire                sleep;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(8),
    .ADDR_WIDTH_B(6),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(128),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("block"),
    .MEMORY_SIZE(32768),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(512),
    .READ_LATENCY_B(2),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(128),
    .WRITE_MODE_B("read_first"),
    .USE_MEM_INIT_MMI(0),
    .WRITE_PROTECT(1)
  ) temp (
    .doutb          (temp_doutb[511:0]), //o
    .addra          (addra[7:0]       ), //i
    .addrb          (addrb[5:0]       ), //i
    .clka           (clk              ), //i
    .clkb           (clk              ), //i
    .dina           (dina[127:0]      ), //i
    .ena            (ena              ), //i
    .enb            (enb              ), //i
    .injectdbiterra (injectdbiterra   ), //i
    .injectsbiterra (injectsbiterra   ), //i
    .regceb         (regceb           ), //i
    .rstb           (rstb             ), //i
    .sleep          (sleep            ), //i
    .wea            (wea              )  //i
  );
  assign injectdbiterra = 1'b0;
  assign injectsbiterra = 1'b0;
  assign regceb = 1'b1;
  assign rstb = 1'b0;
  assign sleep = 1'b0;
  assign doutb = temp_doutb;

endmodule

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

//sdpram replaced by sdpram

module sdpram (
  output     [127:0]  doutb,
  input      [8:0]    addra,
  input      [8:0]    addrb,
  input      [127:0]  dina,
  input               ena,
  input               enb,
  input      [0:0]    wea,
  input               clk
);

  wire       [127:0]  temp_doutb;
  wire                injectdbiterra;
  wire                injectsbiterra;
  wire                regceb;
  wire                rstb;
  wire                sleep;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(128),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("ultra"),
    .MEMORY_SIZE(65536),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(128),
    .READ_LATENCY_B(12),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(128),
    .WRITE_MODE_B("read_first"),
    .USE_MEM_INIT_MMI(0),
    .WRITE_PROTECT(1)
  ) temp (
    .doutb          (temp_doutb[127:0]), //o
    .addra          (addra[8:0]       ), //i
    .addrb          (addrb[8:0]       ), //i
    .clka           (clk              ), //i
    .clkb           (clk              ), //i
    .dina           (dina[127:0]      ), //i
    .ena            (ena              ), //i
    .enb            (enb              ), //i
    .injectdbiterra (injectdbiterra   ), //i
    .injectsbiterra (injectsbiterra   ), //i
    .regceb         (regceb           ), //i
    .rstb           (rstb             ), //i
    .sleep          (sleep            ), //i
    .wea            (wea              )  //i
  );
  assign injectdbiterra = 1'b0;
  assign injectsbiterra = 1'b0;
  assign regceb = 1'b1;
  assign rstb = 1'b0;
  assign sleep = 1'b0;
  assign doutb = temp_doutb;

endmodule

module FeatureConv11Convert (
  input               io_sData_valid,
  output reg          io_sData_ready,
  input      [127:0]  io_sData_payload,
  output              io_mData_mData_0_valid,
  output     [127:0]  io_mData_mData_0_payload,
  output              io_mData_mData_1_valid,
  output     [127:0]  io_mData_mData_1_payload,
  output              io_mData_mData_2_valid,
  output     [127:0]  io_mData_mData_2_payload,
  output              io_mData_mData_3_valid,
  output     [127:0]  io_mData_mData_3_payload,
  output              io_mData_mData_4_valid,
  output     [127:0]  io_mData_mData_4_payload,
  output              io_mData_mData_5_valid,
  output     [127:0]  io_mData_mData_5_payload,
  output              io_mData_mData_6_valid,
  output     [127:0]  io_mData_mData_6_payload,
  output              io_mData_mData_7_valid,
  output     [127:0]  io_mData_mData_7_payload,
  output              io_mData_mData_8_valid,
  output     [127:0]  io_mData_mData_8_payload,
  input               io_mData_ready,
  input      [9:0]    io_rowNumIn,
  input      [9:0]    io_colNumIn,
  input               io_start,
  input      [11:0]   io_channelIn,
  input               clk,
  input               reset,
  input               softReset
);
  localparam FeatureWidthConvertEnum_IDLE = 5'd1;
  localparam FeatureWidthConvertEnum_INIT = 5'd2;
  localparam FeatureWidthConvertEnum_FIFO_READY = 5'd4;
  localparam FeatureWidthConvertEnum_SEND = 5'd8;
  localparam FeatureWidthConvertEnum_END_1 = 5'd16;

  wire       [11:0]   _zz_when_WaCounter_l12_1;
  wire       [7:0]    _zz_when_WaCounter_l12_1_1;
  wire       [9:0]    _zz_when_WaCounter_l12_2;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire                fsm_initEnd;
  wire                fsm_fifoReady;
  wire                fsm_sendEnd;
  wire                fsm_last;
  reg        [4:0]    fsm_currentState;
  reg        [4:0]    fsm_nextState;
  wire                when_WaCounter_l17;
  reg        [2:0]    initCnt_count;
  reg                 initCnt_valid;
  wire                when_WaCounter_l12;
  reg        [7:0]    channelInTimes;
  wire                io_sData_fire;
  reg        [11:0]   channelCnt_count;
  reg                 channelCnt_valid;
  wire                when_WaCounter_l12_1;
  reg        [9:0]    columnCnt_count;
  reg                 columnCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                when_WaCounter_l17_1;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                io_sData_fire_1;
  wire                io_sData_fire_2;
  wire                io_sData_fire_3;
  wire                io_sData_fire_4;
  wire                io_sData_fire_5;
  wire                io_sData_fire_6;
  wire                io_sData_fire_7;
  wire                io_sData_fire_8;
  wire                io_sData_fire_9;
  wire                when_FeatureConv11Convert_l40;
  `ifndef SYNTHESIS
  reg [79:0] fsm_currentState_string;
  reg [79:0] fsm_nextState_string;
  `endif


  assign _zz_when_WaCounter_l12_1_1 = (channelInTimes - 8'h01);
  assign _zz_when_WaCounter_l12_1 = {4'd0, _zz_when_WaCounter_l12_1_1};
  assign _zz_when_WaCounter_l12_2 = (io_colNumIn - 10'h001);
  assign _zz_when_WaCounter_l12_3 = (io_rowNumIn - 10'h001);
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      FeatureWidthConvertEnum_IDLE : fsm_currentState_string = "IDLE      ";
      FeatureWidthConvertEnum_INIT : fsm_currentState_string = "INIT      ";
      FeatureWidthConvertEnum_FIFO_READY : fsm_currentState_string = "FIFO_READY";
      FeatureWidthConvertEnum_SEND : fsm_currentState_string = "SEND      ";
      FeatureWidthConvertEnum_END_1 : fsm_currentState_string = "END_1     ";
      default : fsm_currentState_string = "??????????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      FeatureWidthConvertEnum_IDLE : fsm_nextState_string = "IDLE      ";
      FeatureWidthConvertEnum_INIT : fsm_nextState_string = "INIT      ";
      FeatureWidthConvertEnum_FIFO_READY : fsm_nextState_string = "FIFO_READY";
      FeatureWidthConvertEnum_SEND : fsm_nextState_string = "SEND      ";
      FeatureWidthConvertEnum_END_1 : fsm_nextState_string = "END_1     ";
      default : fsm_nextState_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & FeatureWidthConvertEnum_IDLE) == FeatureWidthConvertEnum_IDLE) : begin
        if(io_start) begin
          fsm_nextState = FeatureWidthConvertEnum_INIT;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_IDLE;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_INIT) == FeatureWidthConvertEnum_INIT) : begin
        if(fsm_initEnd) begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_INIT;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_FIFO_READY) == FeatureWidthConvertEnum_FIFO_READY) : begin
        if(fsm_fifoReady) begin
          fsm_nextState = FeatureWidthConvertEnum_SEND;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_SEND) == FeatureWidthConvertEnum_SEND) : begin
        if(fsm_sendEnd) begin
          fsm_nextState = FeatureWidthConvertEnum_END_1;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_SEND;
        end
      end
      default : begin
        if(fsm_last) begin
          fsm_nextState = FeatureWidthConvertEnum_IDLE;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end
      end
    endcase
  end

  assign when_WaCounter_l17 = ((fsm_currentState & FeatureWidthConvertEnum_INIT) != 5'b00000);
  assign when_WaCounter_l12 = (initCnt_count == 3'b111);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCnt_valid = 1'b1;
    end else begin
      initCnt_valid = 1'b0;
    end
  end

  assign fsm_initEnd = initCnt_valid;
  assign io_sData_fire = (io_sData_valid && io_sData_ready);
  assign when_WaCounter_l12_1 = (channelCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelCnt_valid = 1'b1;
    end else begin
      channelCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l12_2 = (columnCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      columnCnt_valid = 1'b1;
    end else begin
      columnCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_1 = ((fsm_currentState & FeatureWidthConvertEnum_END_1) != 5'b00000);
  assign when_WaCounter_l12_3 = (rowCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
  end

  assign fsm_fifoReady = io_mData_ready;
  assign fsm_sendEnd = (channelCnt_valid && columnCnt_valid);
  assign fsm_last = ((rowCnt_valid && channelCnt_valid) && columnCnt_valid);
  assign io_mData_mData_1_payload = 128'h0;
  assign io_sData_fire_1 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_1_valid = io_sData_fire_1;
  assign io_mData_mData_2_payload = 128'h0;
  assign io_sData_fire_2 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_2_valid = io_sData_fire_2;
  assign io_mData_mData_3_payload = 128'h0;
  assign io_sData_fire_3 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_3_valid = io_sData_fire_3;
  assign io_mData_mData_4_payload = 128'h0;
  assign io_sData_fire_4 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_4_valid = io_sData_fire_4;
  assign io_mData_mData_5_payload = 128'h0;
  assign io_sData_fire_5 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_5_valid = io_sData_fire_5;
  assign io_mData_mData_6_payload = 128'h0;
  assign io_sData_fire_6 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_6_valid = io_sData_fire_6;
  assign io_mData_mData_7_payload = 128'h0;
  assign io_sData_fire_7 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_7_valid = io_sData_fire_7;
  assign io_mData_mData_8_payload = 128'h0;
  assign io_sData_fire_8 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_8_valid = io_sData_fire_8;
  assign io_mData_mData_0_payload = io_sData_payload;
  assign io_sData_fire_9 = (io_sData_valid && io_sData_ready);
  assign io_mData_mData_0_valid = io_sData_fire_9;
  assign when_FeatureConv11Convert_l40 = ((fsm_currentState & FeatureWidthConvertEnum_SEND) != 5'b00000);
  always @(*) begin
    if(when_FeatureConv11Convert_l40) begin
      io_sData_ready = 1'b1;
    end else begin
      io_sData_ready = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      fsm_currentState <= FeatureWidthConvertEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
    end else begin
      if(softReset) begin
      fsm_currentState <= FeatureWidthConvertEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      end else begin
        fsm_currentState <= fsm_nextState;
        if(when_WaCounter_l17) begin
          initCnt_count <= (initCnt_count + 3'b001);
          if(initCnt_valid) begin
            initCnt_count <= 3'b000;
          end
        end
        if(io_sData_fire) begin
          channelCnt_count <= (channelCnt_count + 12'h001);
          if(channelCnt_valid) begin
            channelCnt_count <= 12'h0;
          end
        end
        if(channelCnt_valid) begin
          columnCnt_count <= (columnCnt_count + 10'h001);
          if(columnCnt_valid) begin
            columnCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_1) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    channelInTimes <= (io_channelIn >>> 4);
  end


endmodule

module FeatureWidthConvert (
  input               sData_valid,
  output              sData_ready,
  input      [127:0]  sData_payload,
  output              mData_mData_0_valid,
  output     [127:0]  mData_mData_0_payload,
  output              mData_mData_1_valid,
  output     [127:0]  mData_mData_1_payload,
  output              mData_mData_2_valid,
  output     [127:0]  mData_mData_2_payload,
  output              mData_mData_3_valid,
  output     [127:0]  mData_mData_3_payload,
  output              mData_mData_4_valid,
  output     [127:0]  mData_mData_4_payload,
  output              mData_mData_5_valid,
  output     [127:0]  mData_mData_5_payload,
  output              mData_mData_6_valid,
  output     [127:0]  mData_mData_6_payload,
  output              mData_mData_7_valid,
  output     [127:0]  mData_mData_7_payload,
  output              mData_mData_8_valid,
  output     [127:0]  mData_mData_8_payload,
  input               mData_ready,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input               start,
  input      [11:0]   channelIn,
  input               reset,
  input               clk,
  input               softReset
);
  localparam FeatureWidthConvertEnum_IDLE = 5'd1;
  localparam FeatureWidthConvertEnum_INIT = 5'd2;
  localparam FeatureWidthConvertEnum_FIFO_READY = 5'd4;
  localparam FeatureWidthConvertEnum_SEND = 5'd8;
  localparam FeatureWidthConvertEnum_END_1 = 5'd16;

  reg                 dataCvt_m_axis_tready;
  wire                dataCvt_aresetn;
  wire                dataCvt_s_axis_tready;
  wire                dataCvt_m_axis_tvalid;
  wire       [1023:0] dataCvt_m_axis_tdata;
  wire       [11:0]   _zz_when_WaCounter_l12_1;
  wire       [4:0]    _zz_when_WaCounter_l12_1_1;
  wire       [9:0]    _zz_when_WaCounter_l12_2;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire                fsm_initEnd;
  wire                fsm_fifoReady;
  wire                fsm_sendEnd;
  wire                fsm_last;
  reg        [4:0]    fsm_currentState;
  reg        [4:0]    fsm_nextState;
  wire                when_WaCounter_l17;
  reg        [2:0]    initCnt_count;
  reg                 initCnt_valid;
  wire                when_WaCounter_l12;
  reg        [4:0]    channelInTimes;
  wire                dataCvt_mData_fire;
  reg        [11:0]   channelCnt_count;
  reg                 channelCnt_valid;
  wire                when_WaCounter_l12_1;
  reg        [9:0]    columnCnt_count;
  reg                 columnCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                when_WaCounter_l17_1;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                dataCvt_mData_fire_1;
  wire                dataCvt_mData_fire_2;
  wire                dataCvt_mData_fire_3;
  wire                dataCvt_mData_fire_4;
  wire                dataCvt_mData_fire_5;
  wire                dataCvt_mData_fire_6;
  wire                dataCvt_mData_fire_7;
  wire                dataCvt_mData_fire_8;
  wire                dataCvt_mData_fire_9;
  wire                when_FeatureWidthConvert_l102;
  `ifndef SYNTHESIS
  reg [79:0] fsm_currentState_string;
  reg [79:0] fsm_nextState_string;
  `endif


  assign _zz_when_WaCounter_l12_1_1 = (channelInTimes - 5'h01);
  assign _zz_when_WaCounter_l12_1 = {7'd0, _zz_when_WaCounter_l12_1_1};
  assign _zz_when_WaCounter_l12_2 = (colNumIn - 10'h001);
  assign _zz_when_WaCounter_l12_3 = (rowNumIn - 10'h001);
  conv11DataCvt dataCvt (
    .s_axis_tvalid (sData_valid                 ), //i
    .s_axis_tready (dataCvt_s_axis_tready       ), //o
    .s_axis_tdata  (sData_payload[127:0]        ), //i
    .m_axis_tvalid (dataCvt_m_axis_tvalid       ), //o
    .m_axis_tready (dataCvt_m_axis_tready       ), //i
    .m_axis_tdata  (dataCvt_m_axis_tdata[1023:0]), //o
    .aclk          (clk                         ), //i
    .aresetn       (dataCvt_aresetn             )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      FeatureWidthConvertEnum_IDLE : fsm_currentState_string = "IDLE      ";
      FeatureWidthConvertEnum_INIT : fsm_currentState_string = "INIT      ";
      FeatureWidthConvertEnum_FIFO_READY : fsm_currentState_string = "FIFO_READY";
      FeatureWidthConvertEnum_SEND : fsm_currentState_string = "SEND      ";
      FeatureWidthConvertEnum_END_1 : fsm_currentState_string = "END_1     ";
      default : fsm_currentState_string = "??????????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      FeatureWidthConvertEnum_IDLE : fsm_nextState_string = "IDLE      ";
      FeatureWidthConvertEnum_INIT : fsm_nextState_string = "INIT      ";
      FeatureWidthConvertEnum_FIFO_READY : fsm_nextState_string = "FIFO_READY";
      FeatureWidthConvertEnum_SEND : fsm_nextState_string = "SEND      ";
      FeatureWidthConvertEnum_END_1 : fsm_nextState_string = "END_1     ";
      default : fsm_nextState_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & FeatureWidthConvertEnum_IDLE) == FeatureWidthConvertEnum_IDLE) : begin
        if(start) begin
          fsm_nextState = FeatureWidthConvertEnum_INIT;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_IDLE;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_INIT) == FeatureWidthConvertEnum_INIT) : begin
        if(fsm_initEnd) begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_INIT;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_FIFO_READY) == FeatureWidthConvertEnum_FIFO_READY) : begin
        if(fsm_fifoReady) begin
          fsm_nextState = FeatureWidthConvertEnum_SEND;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end
      end
      (((fsm_currentState) & FeatureWidthConvertEnum_SEND) == FeatureWidthConvertEnum_SEND) : begin
        if(fsm_sendEnd) begin
          fsm_nextState = FeatureWidthConvertEnum_END_1;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_SEND;
        end
      end
      default : begin
        if(fsm_last) begin
          fsm_nextState = FeatureWidthConvertEnum_IDLE;
        end else begin
          fsm_nextState = FeatureWidthConvertEnum_FIFO_READY;
        end
      end
    endcase
  end

  assign when_WaCounter_l17 = ((fsm_currentState & FeatureWidthConvertEnum_INIT) != 5'b00000);
  assign when_WaCounter_l12 = (initCnt_count == 3'b111);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCnt_valid = 1'b1;
    end else begin
      initCnt_valid = 1'b0;
    end
  end

  assign fsm_initEnd = initCnt_valid;
  assign dataCvt_aresetn = (! reset);
  assign dataCvt_mData_fire = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign when_WaCounter_l12_1 = (channelCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelCnt_valid = 1'b1;
    end else begin
      channelCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l12_2 = (columnCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      columnCnt_valid = 1'b1;
    end else begin
      columnCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_1 = ((fsm_currentState & FeatureWidthConvertEnum_END_1) != 5'b00000);
  assign when_WaCounter_l12_3 = (rowCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
  end

  assign fsm_fifoReady = mData_ready;
  assign fsm_sendEnd = (channelCnt_valid && columnCnt_valid);
  assign fsm_last = ((rowCnt_valid && channelCnt_valid) && columnCnt_valid);
  assign sData_ready = dataCvt_s_axis_tready;
  assign mData_mData_0_payload = dataCvt_m_axis_tdata[127 : 0];
  assign dataCvt_mData_fire_1 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_0_valid = dataCvt_mData_fire_1;
  assign mData_mData_1_payload = dataCvt_m_axis_tdata[255 : 128];
  assign dataCvt_mData_fire_2 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_1_valid = dataCvt_mData_fire_2;
  assign mData_mData_2_payload = dataCvt_m_axis_tdata[383 : 256];
  assign dataCvt_mData_fire_3 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_2_valid = dataCvt_mData_fire_3;
  assign mData_mData_3_payload = dataCvt_m_axis_tdata[511 : 384];
  assign dataCvt_mData_fire_4 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_3_valid = dataCvt_mData_fire_4;
  assign mData_mData_4_payload = dataCvt_m_axis_tdata[639 : 512];
  assign dataCvt_mData_fire_5 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_4_valid = dataCvt_mData_fire_5;
  assign mData_mData_5_payload = dataCvt_m_axis_tdata[767 : 640];
  assign dataCvt_mData_fire_6 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_5_valid = dataCvt_mData_fire_6;
  assign mData_mData_6_payload = dataCvt_m_axis_tdata[895 : 768];
  assign dataCvt_mData_fire_7 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_6_valid = dataCvt_mData_fire_7;
  assign mData_mData_7_payload = dataCvt_m_axis_tdata[1023 : 896];
  assign dataCvt_mData_fire_8 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_7_valid = dataCvt_mData_fire_8;
  assign mData_mData_8_payload = 128'h0;
  assign dataCvt_mData_fire_9 = (dataCvt_m_axis_tvalid && dataCvt_m_axis_tready);
  assign mData_mData_8_valid = dataCvt_mData_fire_9;
  assign when_FeatureWidthConvert_l102 = ((fsm_currentState & FeatureWidthConvertEnum_SEND) != 5'b00000);
  always @(*) begin
    if(when_FeatureWidthConvert_l102) begin
      dataCvt_m_axis_tready = 1'b1;
    end else begin
      dataCvt_m_axis_tready = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      fsm_currentState <= FeatureWidthConvertEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
    end else begin
      if(softReset) begin
      fsm_currentState <= FeatureWidthConvertEnum_IDLE;
      initCnt_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      end else begin
        fsm_currentState <= fsm_nextState;
        if(when_WaCounter_l17) begin
          initCnt_count <= (initCnt_count + 3'b001);
          if(initCnt_valid) begin
            initCnt_count <= 3'b000;
          end
        end
        if(dataCvt_mData_fire) begin
          channelCnt_count <= (channelCnt_count + 12'h001);
          if(channelCnt_valid) begin
            channelCnt_count <= 12'h0;
          end
        end
        if(channelCnt_valid) begin
          columnCnt_count <= (columnCnt_count + 10'h001);
          if(columnCnt_valid) begin
            columnCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_1) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    channelInTimes <= (channelIn >>> 7);
  end


endmodule

module FeatureGenerate (
  input               sData_valid,
  output reg          sData_ready,
  input      [127:0]  sData_payload,
  output              mData_mData_0_valid,
  output     [127:0]  mData_mData_0_payload,
  output              mData_mData_1_valid,
  output     [127:0]  mData_mData_1_payload,
  output              mData_mData_2_valid,
  output     [127:0]  mData_mData_2_payload,
  output              mData_mData_3_valid,
  output     [127:0]  mData_mData_3_payload,
  output              mData_mData_4_valid,
  output     [127:0]  mData_mData_4_payload,
  output              mData_mData_5_valid,
  output     [127:0]  mData_mData_5_payload,
  output              mData_mData_6_valid,
  output     [127:0]  mData_mData_6_payload,
  output              mData_mData_7_valid,
  output     [127:0]  mData_mData_7_payload,
  output              mData_mData_8_valid,
  output     [127:0]  mData_mData_8_payload,
  input               mData_ready,
  input      [9:0]    rowNumIn,
  input      [9:0]    colNumIn,
  input               start,
  input      [11:0]   channelIn,
  input               clk,
  input               reset,
  input               softReset
);
  localparam FeatureGenerateEnum_IDLE = 6'd1;
  localparam FeatureGenerateEnum_INIT = 6'd2;
  localparam FeatureGenerateEnum_WAIT_1 = 6'd4;
  localparam FeatureGenerateEnum_FIFO_READY = 6'd8;
  localparam FeatureGenerateEnum_WR = 6'd16;
  localparam FeatureGenerateEnum_END_1 = 6'd32;

  reg        [127:0]  _zz_mem_0_port1;
  reg        [127:0]  _zz_mem_1_port1;
  wire       [17:0]   _zz_when_FeatureGenerate_l129;
  wire       [17:0]   _zz_when_FeatureGenerate_l129_1;
  wire       [127:0]  _zz_mem_0_port;
  wire                _zz_mem_0_port_1;
  wire                _zz_rdData_0;
  wire       [127:0]  _zz_mem_1_port;
  wire                _zz_mem_1_port_1;
  wire                _zz_rdData_1;
  wire       [11:0]   _zz_when_WaCounter_l12_1;
  wire       [7:0]    _zz_when_WaCounter_l12_1_1;
  wire       [9:0]    _zz_when_WaCounter_l12_2;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire       [9:0]    _zz_when_FeatureGenerate_l201;
  wire       [9:0]    _zz_when_FeatureGenerate_l212;
  reg        [7:0]    channelTimes;
  reg        [17:0]   totalCnt;
  wire                fsm_initEnd;
  wire                fsm_waitEnd;
  wire                fsm_wrEnd;
  wire                fsm_endEnd;
  wire                fsm_wait2;
  wire                fsm_fifoReady;
  reg        [5:0]    fsm_currentState;
  reg        [5:0]    fsm_nextState;
  reg        [12:0]   rdAddr;
  wire       [127:0]  wrData_0;
  wire       [127:0]  wrData_1;
  wire       [127:0]  rdData_0;
  wire       [127:0]  rdData_1;
  reg        [12:0]   wrAddr;
  wire                sData_fire;
  wire                when_FeatureGenerate_l129;
  reg        [127:0]  sData_payload_regNext;
  wire                sData_fire_1;
  reg                 sData_fire_1_regNext;
  wire                sData_fire_2;
  reg                 sData_fire_2_regNext;
  wire                when_WaCounter_l17;
  reg        [2:0]    initCount_count;
  reg                 initCount_valid;
  wire                when_WaCounter_l12;
  wire                sData_fire_3;
  reg        [11:0]   channelCnt_count;
  reg                 channelCnt_valid;
  wire                when_WaCounter_l12_1;
  wire                sData_fire_4;
  wire                when_WaCounter_l17_1;
  reg        [9:0]    columnCnt_count;
  reg                 columnCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                when_WaCounter_l17_2;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                when_FeatureGenerate_l191;
  reg                 valid_0;
  reg                 valid_1;
  reg                 valid_2;
  reg                 valid_3;
  reg                 valid_4;
  reg                 valid_5;
  reg                 valid_6;
  reg                 valid_7;
  reg                 valid_8;
  wire                when_FeatureGenerate_l200;
  wire                when_FeatureGenerate_l201;
  wire                when_FeatureGenerate_l212;
  wire                when_FeatureGenerate_l222;
  reg                 valid_0_delay_1;
  reg                 valid_0_delay_2;
  reg                 valid_0_delay_3;
  reg                 valid_3_delay_1;
  reg                 valid_3_delay_2;
  reg                 valid_3_delay_3;
  reg                 valid_6_delay_1;
  reg                 valid_6_delay_2;
  reg                 valid_6_delay_3;
  reg                 valid_1_delay_1;
  reg                 valid_1_delay_2;
  reg                 valid_4_delay_1;
  reg                 valid_4_delay_2;
  reg                 valid_7_delay_1;
  reg                 valid_7_delay_2;
  reg                 valid_2_delay_1;
  reg                 valid_5_delay_1;
  reg                 valid_8_delay_1;
  reg        [127:0]  mData_mData_1_payload_regNext;
  reg        [127:0]  mData_mData_2_payload_regNext;
  reg        [127:0]  rdData_1_regNext;
  reg        [127:0]  mData_mData_4_payload_regNext;
  reg        [127:0]  mData_mData_5_payload_regNext;
  reg        [127:0]  rdData_0_regNext;
  reg        [127:0]  mData_mData_7_payload_regNext;
  reg        [127:0]  mData_mData_8_payload_regNext;
  reg        [127:0]  sData_payload_regNext_1;
  reg        [127:0]  sData_payload_regNext_1_regNext;
  `ifndef SYNTHESIS
  reg [79:0] fsm_currentState_string;
  reg [79:0] fsm_nextState_string;
  `endif

  (* ram_style = "block" *) reg [127:0] mem_0 [0:8191];
  (* ram_style = "block" *) reg [127:0] mem_1 [0:8191];

  assign _zz_when_FeatureGenerate_l129 = {5'd0, rdAddr};
  assign _zz_when_FeatureGenerate_l129_1 = (totalCnt - 18'h00001);
  assign _zz_when_WaCounter_l12_1_1 = (channelTimes - 8'h01);
  assign _zz_when_WaCounter_l12_1 = {4'd0, _zz_when_WaCounter_l12_1_1};
  assign _zz_when_WaCounter_l12_2 = (colNumIn - 10'h001);
  assign _zz_when_WaCounter_l12_3 = (rowNumIn - 10'h001);
  assign _zz_when_FeatureGenerate_l201 = (colNumIn - 10'h002);
  assign _zz_when_FeatureGenerate_l212 = (colNumIn - 10'h001);
  assign _zz_mem_0_port = wrData_0;
  assign _zz_rdData_0 = 1'b1;
  assign _zz_mem_1_port = wrData_1;
  assign _zz_rdData_1 = 1'b1;
  always @(posedge clk) begin
    if(sData_fire_1_regNext) begin
      mem_0[wrAddr] <= _zz_mem_0_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_rdData_0) begin
      _zz_mem_0_port1 <= mem_0[rdAddr];
    end
  end

  always @(posedge clk) begin
    if(sData_fire_2_regNext) begin
      mem_1[wrAddr] <= _zz_mem_1_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_rdData_1) begin
      _zz_mem_1_port1 <= mem_1[rdAddr];
    end
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      FeatureGenerateEnum_IDLE : fsm_currentState_string = "IDLE      ";
      FeatureGenerateEnum_INIT : fsm_currentState_string = "INIT      ";
      FeatureGenerateEnum_WAIT_1 : fsm_currentState_string = "WAIT_1    ";
      FeatureGenerateEnum_FIFO_READY : fsm_currentState_string = "FIFO_READY";
      FeatureGenerateEnum_WR : fsm_currentState_string = "WR        ";
      FeatureGenerateEnum_END_1 : fsm_currentState_string = "END_1     ";
      default : fsm_currentState_string = "??????????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      FeatureGenerateEnum_IDLE : fsm_nextState_string = "IDLE      ";
      FeatureGenerateEnum_INIT : fsm_nextState_string = "INIT      ";
      FeatureGenerateEnum_WAIT_1 : fsm_nextState_string = "WAIT_1    ";
      FeatureGenerateEnum_FIFO_READY : fsm_nextState_string = "FIFO_READY";
      FeatureGenerateEnum_WR : fsm_nextState_string = "WR        ";
      FeatureGenerateEnum_END_1 : fsm_nextState_string = "END_1     ";
      default : fsm_nextState_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & FeatureGenerateEnum_IDLE) == FeatureGenerateEnum_IDLE) : begin
        if(start) begin
          fsm_nextState = FeatureGenerateEnum_INIT;
        end else begin
          fsm_nextState = FeatureGenerateEnum_IDLE;
        end
      end
      (((fsm_currentState) & FeatureGenerateEnum_INIT) == FeatureGenerateEnum_INIT) : begin
        if(fsm_initEnd) begin
          fsm_nextState = FeatureGenerateEnum_WAIT_1;
        end else begin
          fsm_nextState = FeatureGenerateEnum_INIT;
        end
      end
      (((fsm_currentState) & FeatureGenerateEnum_WAIT_1) == FeatureGenerateEnum_WAIT_1) : begin
        if(fsm_waitEnd) begin
          fsm_nextState = FeatureGenerateEnum_END_1;
        end else begin
          fsm_nextState = FeatureGenerateEnum_WAIT_1;
        end
      end
      (((fsm_currentState) & FeatureGenerateEnum_FIFO_READY) == FeatureGenerateEnum_FIFO_READY) : begin
        if(fsm_fifoReady) begin
          fsm_nextState = FeatureGenerateEnum_WR;
        end else begin
          fsm_nextState = FeatureGenerateEnum_FIFO_READY;
        end
      end
      (((fsm_currentState) & FeatureGenerateEnum_WR) == FeatureGenerateEnum_WR) : begin
        if(fsm_wrEnd) begin
          fsm_nextState = FeatureGenerateEnum_END_1;
        end else begin
          fsm_nextState = FeatureGenerateEnum_WR;
        end
      end
      default : begin
        if(fsm_wait2) begin
          fsm_nextState = FeatureGenerateEnum_WAIT_1;
        end else begin
          if(fsm_endEnd) begin
            fsm_nextState = FeatureGenerateEnum_IDLE;
          end else begin
            fsm_nextState = FeatureGenerateEnum_FIFO_READY;
          end
        end
      end
    endcase
  end

  assign fsm_fifoReady = mData_ready;
  assign sData_fire = (sData_valid && sData_ready);
  assign when_FeatureGenerate_l129 = (_zz_when_FeatureGenerate_l129 == _zz_when_FeatureGenerate_l129_1);
  assign wrData_0 = sData_payload_regNext;
  assign wrData_1 = rdData_0;
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign rdData_0 = _zz_mem_0_port1;
  assign sData_fire_2 = (sData_valid && sData_ready);
  assign rdData_1 = _zz_mem_1_port1;
  assign when_WaCounter_l17 = ((fsm_currentState & FeatureGenerateEnum_INIT) != 6'b000000);
  assign when_WaCounter_l12 = (initCount_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCount_valid = 1'b1;
    end else begin
      initCount_valid = 1'b0;
    end
  end

  assign fsm_initEnd = initCount_valid;
  assign sData_fire_3 = (sData_valid && sData_ready);
  assign when_WaCounter_l12_1 = (channelCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelCnt_valid = 1'b1;
    end else begin
      channelCnt_valid = 1'b0;
    end
  end

  assign sData_fire_4 = (sData_valid && sData_ready);
  assign when_WaCounter_l17_1 = (channelCnt_valid && sData_fire_4);
  assign when_WaCounter_l12_2 = (columnCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      columnCnt_valid = 1'b1;
    end else begin
      columnCnt_valid = 1'b0;
    end
  end

  assign when_WaCounter_l17_2 = ((fsm_currentState & FeatureGenerateEnum_END_1) != 6'b000000);
  assign when_WaCounter_l12_3 = (rowCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
  end

  assign fsm_waitEnd = (channelCnt_valid && columnCnt_valid);
  assign fsm_wait2 = (rowCnt_count < 10'h001);
  assign fsm_wrEnd = (channelCnt_valid && columnCnt_valid);
  assign fsm_endEnd = rowCnt_valid;
  assign when_FeatureGenerate_l191 = (((fsm_currentState & FeatureGenerateEnum_WAIT_1) != 6'b000000) || ((fsm_currentState & FeatureGenerateEnum_WR) != 6'b000000));
  always @(*) begin
    if(when_FeatureGenerate_l191) begin
      sData_ready = 1'b1;
    end else begin
      sData_ready = 1'b0;
    end
  end

  assign when_FeatureGenerate_l200 = ((fsm_currentState & FeatureGenerateEnum_WR) != 6'b000000);
  assign when_FeatureGenerate_l201 = (columnCnt_count < _zz_when_FeatureGenerate_l201);
  assign when_FeatureGenerate_l212 = ((10'h0 < columnCnt_count) && (columnCnt_count < _zz_when_FeatureGenerate_l212));
  assign when_FeatureGenerate_l222 = ((10'h001 < columnCnt_count) && (columnCnt_count < colNumIn));
  assign mData_mData_0_valid = valid_0_delay_3;
  assign mData_mData_3_valid = valid_3_delay_3;
  assign mData_mData_6_valid = valid_6_delay_3;
  assign mData_mData_1_valid = valid_1_delay_2;
  assign mData_mData_4_valid = valid_4_delay_2;
  assign mData_mData_7_valid = valid_7_delay_2;
  assign mData_mData_2_valid = valid_2_delay_1;
  assign mData_mData_5_valid = valid_5_delay_1;
  assign mData_mData_8_valid = valid_8_delay_1;
  assign mData_mData_0_payload = mData_mData_1_payload_regNext;
  assign mData_mData_1_payload = mData_mData_2_payload_regNext;
  assign mData_mData_2_payload = rdData_1_regNext;
  assign mData_mData_3_payload = mData_mData_4_payload_regNext;
  assign mData_mData_4_payload = mData_mData_5_payload_regNext;
  assign mData_mData_5_payload = rdData_0_regNext;
  assign mData_mData_6_payload = mData_mData_7_payload_regNext;
  assign mData_mData_7_payload = mData_mData_8_payload_regNext;
  assign mData_mData_8_payload = sData_payload_regNext_1_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      channelTimes <= 8'h0;
      fsm_currentState <= FeatureGenerateEnum_IDLE;
      rdAddr <= 13'h0;
      initCount_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      valid_0 <= 1'b0;
      valid_1 <= 1'b0;
      valid_2 <= 1'b0;
      valid_3 <= 1'b0;
      valid_4 <= 1'b0;
      valid_5 <= 1'b0;
      valid_6 <= 1'b0;
      valid_7 <= 1'b0;
      valid_8 <= 1'b0;
    end else begin
      if(softReset) begin
      channelTimes <= 8'h0;
      fsm_currentState <= FeatureGenerateEnum_IDLE;
      rdAddr <= 13'h0;
      initCount_count <= 3'b000;
      channelCnt_count <= 12'h0;
      columnCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      valid_0 <= 1'b0;
      valid_1 <= 1'b0;
      valid_2 <= 1'b0;
      valid_3 <= 1'b0;
      valid_4 <= 1'b0;
      valid_5 <= 1'b0;
      valid_6 <= 1'b0;
      valid_7 <= 1'b0;
      valid_8 <= 1'b0;
      end else begin
        channelTimes <= (channelIn >>> 4);
        fsm_currentState <= fsm_nextState;
        if(sData_fire) begin
          if(when_FeatureGenerate_l129) begin
            rdAddr <= 13'h0;
          end else begin
            rdAddr <= (rdAddr + 13'h0001);
          end
        end
        if(when_WaCounter_l17) begin
          initCount_count <= (initCount_count + 3'b001);
          if(initCount_valid) begin
            initCount_count <= 3'b000;
          end
        end
        if(sData_fire_3) begin
          channelCnt_count <= (channelCnt_count + 12'h001);
          if(channelCnt_valid) begin
            channelCnt_count <= 12'h0;
          end
        end
        if(when_WaCounter_l17_1) begin
          columnCnt_count <= (columnCnt_count + 10'h001);
          if(columnCnt_valid) begin
            columnCnt_count <= 10'h0;
          end
        end
        if(when_WaCounter_l17_2) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
        if(when_FeatureGenerate_l200) begin
          if(when_FeatureGenerate_l201) begin
            valid_0 <= 1'b1;
            valid_3 <= 1'b1;
            valid_6 <= 1'b1;
          end else begin
            valid_0 <= 1'b0;
            valid_3 <= 1'b0;
            valid_6 <= 1'b0;
          end
          if(when_FeatureGenerate_l212) begin
            valid_1 <= 1'b1;
            valid_4 <= 1'b1;
            valid_7 <= 1'b1;
          end else begin
            valid_1 <= 1'b0;
            valid_4 <= 1'b0;
            valid_7 <= 1'b0;
          end
          if(when_FeatureGenerate_l222) begin
            valid_2 <= 1'b1;
            valid_5 <= 1'b1;
            valid_8 <= 1'b1;
          end else begin
            valid_2 <= 1'b0;
            valid_5 <= 1'b0;
            valid_8 <= 1'b0;
          end
        end else begin
          valid_0 <= 1'b0;
          valid_1 <= 1'b0;
          valid_2 <= 1'b0;
          valid_3 <= 1'b0;
          valid_4 <= 1'b0;
          valid_5 <= 1'b0;
          valid_6 <= 1'b0;
          valid_7 <= 1'b0;
          valid_8 <= 1'b0;
        end
      end
    end
  end

  always @(posedge clk) begin
    totalCnt <= (channelTimes * colNumIn);
    wrAddr <= rdAddr;
    sData_payload_regNext <= sData_payload;
    sData_fire_1_regNext <= sData_fire_1;
    sData_fire_2_regNext <= sData_fire_2;
    valid_0_delay_1 <= valid_0;
    valid_0_delay_2 <= valid_0_delay_1;
    valid_0_delay_3 <= valid_0_delay_2;
    valid_3_delay_1 <= valid_3;
    valid_3_delay_2 <= valid_3_delay_1;
    valid_3_delay_3 <= valid_3_delay_2;
    valid_6_delay_1 <= valid_6;
    valid_6_delay_2 <= valid_6_delay_1;
    valid_6_delay_3 <= valid_6_delay_2;
    valid_1_delay_1 <= valid_1;
    valid_1_delay_2 <= valid_1_delay_1;
    valid_4_delay_1 <= valid_4;
    valid_4_delay_2 <= valid_4_delay_1;
    valid_7_delay_1 <= valid_7;
    valid_7_delay_2 <= valid_7_delay_1;
    valid_2_delay_1 <= valid_2;
    valid_5_delay_1 <= valid_5;
    valid_8_delay_1 <= valid_8;
    mData_mData_1_payload_regNext <= mData_mData_1_payload;
    mData_mData_2_payload_regNext <= mData_mData_2_payload;
    rdData_1_regNext <= rdData_1;
    mData_mData_4_payload_regNext <= mData_mData_4_payload;
    mData_mData_5_payload_regNext <= mData_mData_5_payload;
    rdData_0_regNext <= rdData_0;
    mData_mData_7_payload_regNext <= mData_mData_7_payload;
    mData_mData_8_payload_regNext <= mData_mData_8_payload;
    sData_payload_regNext_1 <= sData_payload;
    sData_payload_regNext_1_regNext <= sData_payload_regNext_1;
  end


endmodule

module Padding (
  input               sData_valid,
  output              sData_ready,
  input      [127:0]  sData_payload,
  output              mData_valid,
  input               mData_ready,
  output     [127:0]  mData_payload,
  input               enPadding,
  input      [11:0]   channelIn,
  input               start,
  input      [9:0]    rowNumIn,
  output reg [9:0]    rowNumOut,
  input      [9:0]    colNumIn,
  output reg [9:0]    colNumOut,
  input      [7:0]    zeroDara,
  input      [0:0]    zeroNum,
  input               clk,
  input               reset,
  input               softReset
);
  localparam PaddingEnum_IDLE = 7'd1;
  localparam PaddingEnum_INIT = 7'd2;
  localparam PaddingEnum_UPDOWN = 7'd4;
  localparam PaddingEnum_LEFT = 7'd8;
  localparam PaddingEnum_CENTER = 7'd16;
  localparam PaddingEnum_RIGHT = 7'd32;
  localparam PaddingEnum_END_1 = 7'd64;

  reg                 fifo_push_valid;
  reg        [127:0]  fifo_push_payload;
  wire                fifo_push_ready;
  wire                fifo_pop_valid;
  wire       [127:0]  fifo_pop_payload;
  wire       [9:0]    _zz_rowNumOut;
  wire       [1:0]    _zz_rowNumOut_1;
  wire       [9:0]    _zz_colNumOut;
  wire       [1:0]    _zz_colNumOut_1;
  wire       [11:0]   _zz_when_WaCounter_l12_1;
  wire       [7:0]    _zz_when_WaCounter_l12_1_1;
  wire       [9:0]    _zz_when_WaCounter_l12_2;
  wire       [9:0]    _zz_when_WaCounter_l12_3;
  wire       [9:0]    _zz_when_Padding_l179_1;
  wire       [0:0]    _zz_when_Padding_l179_1_1;
  wire       [9:0]    _zz_when_Padding_l179_2;
  wire       [9:0]    _zz_when_Padding_l179_3;
  wire       [9:0]    _zz_when_Padding_l179_4;
  wire       [9:0]    _zz_when_Padding_l179_4_1;
  wire       [9:0]    _zz_when_Padding_l179_4_2;
  wire       [9:0]    _zz_when_Padding_l179_5;
  wire       [9:0]    _zz_when_Padding_l179_5_1;
  wire       [9:0]    _zz_when_Padding_l179_5_2;
  wire       [9:0]    _zz_when_Padding_l179_6;
  wire       [9:0]    _zz_when_Padding_l179_6_1;
  wire       [9:0]    _zz_when_Padding_l179_6_2;
  wire       [9:0]    _zz_when_Padding_l179_6_3;
  reg        [7:0]    channelTimes;
  wire                fsm_initEnd;
  reg                 fsm_leftEnd;
  reg                 fsm_rightEnd;
  reg                 fsm_upDownEnd;
  reg                 fsm_centerEnd;
  reg                 fsm_endEnd;
  wire                fsm_enPadding;
  reg                 fsm_enUpDown;
  reg        [6:0]    fsm_currentState;
  reg        [6:0]    fsm_nextState;
  reg                 initEn;
  wire                when_Padding_l186;
  wire                when_Padding_l186_1;
  reg        [4:0]    initCount_count;
  reg                 initCount_valid;
  wire                when_WaCounter_l12;
  wire                when_Padding_l190;
  reg                 zeroValid;
  wire                when_Padding_l197;
  wire       [7:0]    _zz_push_payload;
  wire                fifo_push_fire;
  reg        [11:0]   channelCnt_count;
  reg                 channelCnt_valid;
  wire                when_WaCounter_l12_1;
  wire                when_Padding_l213;
  wire                fifo_push_fire_1;
  wire                when_WaCounter_l17;
  reg        [9:0]    colCnt_count;
  reg                 colCnt_valid;
  wire                when_WaCounter_l12_2;
  wire                when_Padding_l220;
  wire                when_WaCounter_l17_1;
  reg        [9:0]    rowCnt_count;
  reg                 rowCnt_valid;
  wire                when_WaCounter_l12_3;
  wire                when_Padding_l227;
  wire                when_Padding_l179;
  wire                fifo_push_fire_2;
  wire                when_Padding_l179_1;
  wire                fifo_push_fire_3;
  wire                when_Padding_l179_2;
  wire                when_Padding_l179_3;
  wire                fifo_push_fire_4;
  wire                when_Padding_l179_4;
  wire                fifo_push_fire_5;
  wire                when_Padding_l179_5;
  wire                when_Padding_l179_6;
  `ifndef SYNTHESIS
  reg [47:0] fsm_currentState_string;
  reg [47:0] fsm_nextState_string;
  `endif


  assign _zz_rowNumOut_1 = ({1'd0,zeroNum} <<< 1);
  assign _zz_rowNumOut = {8'd0, _zz_rowNumOut_1};
  assign _zz_colNumOut_1 = ({1'd0,zeroNum} <<< 1);
  assign _zz_colNumOut = {8'd0, _zz_colNumOut_1};
  assign _zz_when_WaCounter_l12_1_1 = (channelTimes - 8'h01);
  assign _zz_when_WaCounter_l12_1 = {4'd0, _zz_when_WaCounter_l12_1_1};
  assign _zz_when_WaCounter_l12_2 = (colNumOut - 10'h001);
  assign _zz_when_WaCounter_l12_3 = (rowNumOut - 10'h001);
  assign _zz_when_Padding_l179_1_1 = (zeroNum - 1'b1);
  assign _zz_when_Padding_l179_1 = {9'd0, _zz_when_Padding_l179_1_1};
  assign _zz_when_Padding_l179_2 = (colNumOut - 10'h001);
  assign _zz_when_Padding_l179_3 = (rowNumOut - 10'h001);
  assign _zz_when_Padding_l179_4 = (_zz_when_Padding_l179_4_1 - 10'h001);
  assign _zz_when_Padding_l179_4_1 = (colNumOut - _zz_when_Padding_l179_4_2);
  assign _zz_when_Padding_l179_4_2 = {9'd0, zeroNum};
  assign _zz_when_Padding_l179_5 = (_zz_when_Padding_l179_5_1 - 10'h001);
  assign _zz_when_Padding_l179_5_1 = (colNumOut - _zz_when_Padding_l179_5_2);
  assign _zz_when_Padding_l179_5_2 = {9'd0, zeroNum};
  assign _zz_when_Padding_l179_6 = {9'd0, zeroNum};
  assign _zz_when_Padding_l179_6_1 = (_zz_when_Padding_l179_6_2 - 10'h001);
  assign _zz_when_Padding_l179_6_2 = (rowNumOut - _zz_when_Padding_l179_6_3);
  assign _zz_when_Padding_l179_6_3 = {9'd0, zeroNum};
  WaStreamFifo fifo (
    .push_valid   (fifo_push_valid         ), //i
    .push_ready   (fifo_push_ready         ), //o
    .push_payload (fifo_push_payload[127:0]), //i
    .pop_valid    (fifo_pop_valid          ), //o
    .pop_ready    (mData_ready             ), //i
    .pop_payload  (fifo_pop_payload[127:0] ), //o
    .flush        (1'b0                    ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   ), //i
    .softReset    (softReset               )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_currentState)
      PaddingEnum_IDLE : fsm_currentState_string = "IDLE  ";
      PaddingEnum_INIT : fsm_currentState_string = "INIT  ";
      PaddingEnum_UPDOWN : fsm_currentState_string = "UPDOWN";
      PaddingEnum_LEFT : fsm_currentState_string = "LEFT  ";
      PaddingEnum_CENTER : fsm_currentState_string = "CENTER";
      PaddingEnum_RIGHT : fsm_currentState_string = "RIGHT ";
      PaddingEnum_END_1 : fsm_currentState_string = "END_1 ";
      default : fsm_currentState_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_nextState)
      PaddingEnum_IDLE : fsm_nextState_string = "IDLE  ";
      PaddingEnum_INIT : fsm_nextState_string = "INIT  ";
      PaddingEnum_UPDOWN : fsm_nextState_string = "UPDOWN";
      PaddingEnum_LEFT : fsm_nextState_string = "LEFT  ";
      PaddingEnum_CENTER : fsm_nextState_string = "CENTER";
      PaddingEnum_RIGHT : fsm_nextState_string = "RIGHT ";
      PaddingEnum_END_1 : fsm_nextState_string = "END_1 ";
      default : fsm_nextState_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    if(enPadding) begin
      rowNumOut = (_zz_rowNumOut + rowNumIn);
    end else begin
      rowNumOut = rowNumIn;
    end
  end

  always @(*) begin
    if(enPadding) begin
      colNumOut = (_zz_colNumOut + colNumIn);
    end else begin
      colNumOut = colNumIn;
    end
  end

  assign mData_valid = fifo_pop_valid;
  assign mData_payload = fifo_pop_payload;
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_currentState) & PaddingEnum_IDLE) == PaddingEnum_IDLE) : begin
        if(start) begin
          fsm_nextState = PaddingEnum_INIT;
        end else begin
          fsm_nextState = PaddingEnum_IDLE;
        end
      end
      (((fsm_currentState) & PaddingEnum_INIT) == PaddingEnum_INIT) : begin
        if(fsm_initEnd) begin
          if(fsm_enPadding) begin
            fsm_nextState = PaddingEnum_LEFT;
          end else begin
            fsm_nextState = PaddingEnum_CENTER;
          end
        end else begin
          fsm_nextState = PaddingEnum_INIT;
        end
      end
      (((fsm_currentState) & PaddingEnum_UPDOWN) == PaddingEnum_UPDOWN) : begin
        if(fsm_upDownEnd) begin
          fsm_nextState = PaddingEnum_RIGHT;
        end else begin
          fsm_nextState = PaddingEnum_UPDOWN;
        end
      end
      (((fsm_currentState) & PaddingEnum_LEFT) == PaddingEnum_LEFT) : begin
        if(fsm_leftEnd) begin
          if(fsm_enUpDown) begin
            fsm_nextState = PaddingEnum_UPDOWN;
          end else begin
            fsm_nextState = PaddingEnum_CENTER;
          end
        end else begin
          fsm_nextState = PaddingEnum_LEFT;
        end
      end
      (((fsm_currentState) & PaddingEnum_CENTER) == PaddingEnum_CENTER) : begin
        if(fsm_centerEnd) begin
          if(fsm_enPadding) begin
            fsm_nextState = PaddingEnum_RIGHT;
          end else begin
            fsm_nextState = PaddingEnum_END_1;
          end
        end else begin
          fsm_nextState = PaddingEnum_CENTER;
        end
      end
      (((fsm_currentState) & PaddingEnum_RIGHT) == PaddingEnum_RIGHT) : begin
        if(fsm_rightEnd) begin
          fsm_nextState = PaddingEnum_END_1;
        end else begin
          fsm_nextState = PaddingEnum_RIGHT;
        end
      end
      default : begin
        if(fsm_endEnd) begin
          fsm_nextState = PaddingEnum_IDLE;
        end else begin
          if(fsm_enPadding) begin
            fsm_nextState = PaddingEnum_LEFT;
          end else begin
            fsm_nextState = PaddingEnum_CENTER;
          end
        end
      end
    endcase
  end

  assign fsm_enPadding = enPadding;
  assign sData_ready = (fifo_push_ready && ((fsm_currentState & PaddingEnum_CENTER) != 7'b0000000));
  assign when_Padding_l186 = ((fsm_currentState & PaddingEnum_INIT) != 7'b0000000);
  assign when_Padding_l186_1 = ((fsm_nextState & PaddingEnum_INIT) == 7'b0000000);
  assign when_WaCounter_l12 = (initCount_count == 5'h08);
  always @(*) begin
    if(when_WaCounter_l12) begin
      initCount_valid = 1'b1;
    end else begin
      initCount_valid = 1'b0;
    end
    if(when_Padding_l190) begin
      initCount_valid = 1'b0;
    end
  end

  assign when_Padding_l190 = ((fsm_currentState & PaddingEnum_IDLE) != 7'b0000000);
  assign fsm_initEnd = initCount_valid;
  assign when_Padding_l197 = ((fsm_currentState & PaddingEnum_CENTER) != 7'b0000000);
  always @(*) begin
    if(when_Padding_l197) begin
      fifo_push_valid = sData_valid;
    end else begin
      fifo_push_valid = zeroValid;
    end
  end

  always @(*) begin
    if(when_Padding_l197) begin
      fifo_push_payload = sData_payload;
    end else begin
      fifo_push_payload[7 : 0] = _zz_push_payload;
      fifo_push_payload[15 : 8] = _zz_push_payload;
      fifo_push_payload[23 : 16] = _zz_push_payload;
      fifo_push_payload[31 : 24] = _zz_push_payload;
      fifo_push_payload[39 : 32] = _zz_push_payload;
      fifo_push_payload[47 : 40] = _zz_push_payload;
      fifo_push_payload[55 : 48] = _zz_push_payload;
      fifo_push_payload[63 : 56] = _zz_push_payload;
      fifo_push_payload[71 : 64] = _zz_push_payload;
      fifo_push_payload[79 : 72] = _zz_push_payload;
      fifo_push_payload[87 : 80] = _zz_push_payload;
      fifo_push_payload[95 : 88] = _zz_push_payload;
      fifo_push_payload[103 : 96] = _zz_push_payload;
      fifo_push_payload[111 : 104] = _zz_push_payload;
      fifo_push_payload[119 : 112] = _zz_push_payload;
      fifo_push_payload[127 : 120] = _zz_push_payload;
    end
  end

  assign _zz_push_payload = zeroDara;
  assign fifo_push_fire = (fifo_push_valid && fifo_push_ready);
  assign when_WaCounter_l12_1 = (channelCnt_count == _zz_when_WaCounter_l12_1);
  always @(*) begin
    if(when_WaCounter_l12_1) begin
      channelCnt_valid = 1'b1;
    end else begin
      channelCnt_valid = 1'b0;
    end
    if(when_Padding_l213) begin
      channelCnt_valid = 1'b0;
    end
  end

  assign when_Padding_l213 = ((fsm_currentState & PaddingEnum_IDLE) != 7'b0000000);
  assign fifo_push_fire_1 = (fifo_push_valid && fifo_push_ready);
  assign when_WaCounter_l17 = (channelCnt_valid && fifo_push_fire_1);
  assign when_WaCounter_l12_2 = (colCnt_count == _zz_when_WaCounter_l12_2);
  always @(*) begin
    if(when_WaCounter_l12_2) begin
      colCnt_valid = 1'b1;
    end else begin
      colCnt_valid = 1'b0;
    end
    if(when_Padding_l220) begin
      colCnt_valid = 1'b0;
    end
  end

  assign when_Padding_l220 = ((fsm_currentState & PaddingEnum_IDLE) != 7'b0000000);
  assign when_WaCounter_l17_1 = ((fsm_nextState & PaddingEnum_END_1) != 7'b0000000);
  assign when_WaCounter_l12_3 = (rowCnt_count == _zz_when_WaCounter_l12_3);
  always @(*) begin
    if(when_WaCounter_l12_3) begin
      rowCnt_valid = 1'b1;
    end else begin
      rowCnt_valid = 1'b0;
    end
    if(when_Padding_l227) begin
      rowCnt_valid = 1'b0;
    end
  end

  assign when_Padding_l227 = ((fsm_currentState & PaddingEnum_IDLE) != 7'b0000000);
  assign when_Padding_l179 = ((((fsm_currentState & PaddingEnum_LEFT) != 7'b0000000) || ((fsm_currentState & PaddingEnum_RIGHT) != 7'b0000000)) || ((fsm_currentState & PaddingEnum_UPDOWN) != 7'b0000000));
  always @(*) begin
    if(when_Padding_l179) begin
      zeroValid = 1'b1;
    end else begin
      zeroValid = 1'b0;
    end
  end

  assign fifo_push_fire_2 = (fifo_push_valid && fifo_push_ready);
  assign when_Padding_l179_1 = (((colCnt_count == _zz_when_Padding_l179_1) && channelCnt_valid) && fifo_push_fire_2);
  always @(*) begin
    if(when_Padding_l179_1) begin
      fsm_leftEnd = 1'b1;
    end else begin
      fsm_leftEnd = 1'b0;
    end
  end

  assign fifo_push_fire_3 = (fifo_push_valid && fifo_push_ready);
  assign when_Padding_l179_2 = (((colCnt_count == _zz_when_Padding_l179_2) && channelCnt_valid) && fifo_push_fire_3);
  always @(*) begin
    if(when_Padding_l179_2) begin
      fsm_rightEnd = 1'b1;
    end else begin
      fsm_rightEnd = 1'b0;
    end
  end

  assign when_Padding_l179_3 = (rowCnt_count == _zz_when_Padding_l179_3);
  assign fifo_push_fire_4 = (fifo_push_valid && fifo_push_ready);
  assign when_Padding_l179_4 = (((colCnt_count == _zz_when_Padding_l179_4) && channelCnt_valid) && fifo_push_fire_4);
  always @(*) begin
    if(when_Padding_l179_4) begin
      fsm_upDownEnd = 1'b1;
    end else begin
      fsm_upDownEnd = 1'b0;
    end
  end

  assign fifo_push_fire_5 = (fifo_push_valid && fifo_push_ready);
  assign when_Padding_l179_5 = (((colCnt_count == _zz_when_Padding_l179_5) && channelCnt_valid) && fifo_push_fire_5);
  always @(*) begin
    if(when_Padding_l179_5) begin
      fsm_centerEnd = 1'b1;
    end else begin
      fsm_centerEnd = 1'b0;
    end
  end

  assign when_Padding_l179_6 = ((rowCnt_count < _zz_when_Padding_l179_6) || (_zz_when_Padding_l179_6_1 < rowCnt_count));
  always @(*) begin
    if(when_Padding_l179_6) begin
      fsm_enUpDown = 1'b1;
    end else begin
      fsm_enUpDown = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      channelTimes <= 8'h0;
      fsm_currentState <= PaddingEnum_IDLE;
      initEn <= 1'b0;
      initCount_count <= 5'h0;
      channelCnt_count <= 12'h0;
      colCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
    end else begin
      if(softReset) begin
      channelTimes <= 8'h0;
      fsm_currentState <= PaddingEnum_IDLE;
      initEn <= 1'b0;
      initCount_count <= 5'h0;
      channelCnt_count <= 12'h0;
      colCnt_count <= 10'h0;
      rowCnt_count <= 10'h0;
      end else begin
        channelTimes <= (channelIn >>> 4);
        fsm_currentState <= fsm_nextState;
        if(when_Padding_l186) begin
          initEn <= 1'b1;
        end
        if(when_Padding_l186_1) begin
          initEn <= 1'b0;
        end
        if(initEn) begin
          initCount_count <= (initCount_count + 5'h01);
          if(initCount_valid) begin
            initCount_count <= 5'h0;
          end
        end
        if(when_Padding_l190) begin
          initCount_count <= 5'h0;
        end
        if(fifo_push_fire) begin
          channelCnt_count <= (channelCnt_count + 12'h001);
          if(channelCnt_valid) begin
            channelCnt_count <= 12'h0;
          end
        end
        if(when_Padding_l213) begin
          channelCnt_count <= 12'h0;
        end
        if(when_WaCounter_l17) begin
          colCnt_count <= (colCnt_count + 10'h001);
          if(colCnt_valid) begin
            colCnt_count <= 10'h0;
          end
        end
        if(when_Padding_l220) begin
          colCnt_count <= 10'h0;
        end
        if(when_WaCounter_l17_1) begin
          rowCnt_count <= (rowCnt_count + 10'h001);
          if(rowCnt_valid) begin
            rowCnt_count <= 10'h0;
          end
        end
        if(when_Padding_l227) begin
          rowCnt_count <= 10'h0;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(when_Padding_l179_3) begin
      fsm_endEnd <= 1'b1;
    end else begin
      fsm_endEnd <= 1'b0;
    end
  end


endmodule

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [127:0]  io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [127:0]  io_pop_payload,
  input               io_flush,
  output     [14:0]   io_availability,
  input               clk,
  input               reset,
  input               softReset
);

  reg        [127:0]  _zz_logic_ram_port0;
  wire       [13:0]   _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [13:0]   _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [127:0]  _zz_logic_ram_port_1;
  wire       [13:0]   _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [13:0]   logic_pushPtr_valueNext;
  reg        [13:0]   logic_pushPtr_value;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [13:0]   logic_popPtr_valueNext;
  reg        [13:0]   logic_popPtr_value;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1075;
  reg [127:0] logic_ram [0:16383];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {13'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {13'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 14'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 14'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 14'h0;
      logic_popPtr_value <= 14'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      if(softReset) begin
      logic_pushPtr_value <= 14'h0;
      logic_popPtr_value <= 14'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
      end else begin
        logic_pushPtr_value <= logic_pushPtr_valueNext;
        logic_popPtr_value <= logic_popPtr_valueNext;
        _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
        if(when_Stream_l1075) begin
          logic_risingOccupancy <= logic_pushing;
        end
        if(io_flush) begin
          logic_risingOccupancy <= 1'b0;
        end
      end
    end
  end


endmodule

module WaStreamFifo (
  input               push_valid,
  output              push_ready,
  input      [127:0]  push_payload,
  output              pop_valid,
  input               pop_ready,
  output     [127:0]  pop_payload,
  input               flush,
  input               clk,
  input               reset,
  input               softReset
);

  reg        [127:0]  _zz_logic_ram_port0;
  wire       [2:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [2:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_pop_payload;
  wire       [127:0]  _zz_logic_ram_port_1;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [2:0]    logic_pushPtr_valueNext;
  reg        [2:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [2:0]    logic_popPtr_valueNext;
  reg        [2:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_pop_valid;
  wire                when_Stream_l1075;
  reg [127:0] logic_ram [0:4];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {2'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {2'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = push_payload;
  always @(posedge clk) begin
    if(_zz_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 3'b100);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    if(logic_pushPtr_willOverflow) begin
      logic_pushPtr_valueNext = 3'b000;
    end else begin
      logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    end
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 3'b000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 3'b100);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    if(logic_popPtr_willOverflow) begin
      logic_popPtr_valueNext = 3'b000;
    end else begin
      logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    end
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 3'b000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (push_valid && push_ready);
  assign logic_popping = (pop_valid && pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign push_ready = (! logic_full);
  assign pop_valid = ((! logic_empty) && (! (_zz_pop_valid && (! logic_full))));
  assign pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 3'b000;
      logic_popPtr_value <= 3'b000;
      logic_risingOccupancy <= 1'b0;
      _zz_pop_valid <= 1'b0;
    end else begin
      if(softReset) begin
      logic_pushPtr_value <= 3'b000;
      logic_popPtr_value <= 3'b000;
      logic_risingOccupancy <= 1'b0;
      _zz_pop_valid <= 1'b0;
      end else begin
        logic_pushPtr_value <= logic_pushPtr_valueNext;
        logic_popPtr_value <= logic_popPtr_valueNext;
        _zz_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
        if(when_Stream_l1075) begin
          logic_risingOccupancy <= logic_pushing;
        end
        if(flush) begin
          logic_risingOccupancy <= 1'b0;
        end
      end
    end
  end


endmodule

module DSP (
              input             [7:0] a       ,
              input             [7:0] d       ,
              input             [7:0] b       ,
              output   reg      [31:0] p      ,
              input             CLK

          );

          wire  signed       [7:0]   ain;
          assign ain = $signed(a);
          wire  signed       [24:0]  din;
          wire [33:0] pout;
          wire [15:0] a1;
          wire [15:0] a2;
          assign a1 = pout[15:0];
          assign a2 = pout[31:16];
          always@(*)begin
               if(a1[15])begin
                   p[15:0] = a1;
                   p[31:16] = a2+1;
               end else begin
                   p[15:0] = a1;
                   p[31:16] = a2;
               end
          end
          assign din =  $signed({d,16'd0});
          mulWeight mulWeight_inst (
            .CLK(CLK),  // input wire CLK
            .A(ain),      // input wire [7 : 0] A
            .B({1'b0,b}),      // input wire [8 : 0] B
            .D(din),      // input wire [24 : 0] D
            .P(pout)      // output wire [33 : 0] P
          );

endmodule
      
